* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py

.SUBCKT s_equivalent p1 p2 p3 p4 p5 p6 p7 p8 p9 p10 p11 p12 p13 p14 p15 p16

* Port network for port 1
R_ref_1 p1 a1 50.0
H_b_1 a1 0 V_c_1 14.142135623730951
* Differential incident wave a sources for transfer from port 1
H_p_1 nt_p_1 nts_p_1 H_b_1 3.5355339059327378
E_p_1 nts_p_1 0 p1 0 0.07071067811865475
E_n_1 0 nt_n_1 nt_p_1 0 1
* Current sensor on center node for transfer to port 1
V_c_1 nt_c_1 0 0
* Transfer network from port 1 to port 1
R1_1 nt_n_1 nt_c_1 3.055402905354145
X1 nt_n_1 nt_c_1 rl_admittance res=1.565082328677509 ind=1.3504716875466727e-07
X2 nt_n_1 nt_c_1 rl_admittance res=20.133594041960766 ind=7.695994849647124e-06
X3 nt_p_1 nt_c_1 rl_admittance res=40.50019708855462 ind=3.3998907307601685e-05
X4 nt_n_1 nt_c_1 rl_admittance res=10.606969280684247 ind=0.0003605354379150948
X5 nt_n_1 nt_c_1 rl_admittance res=1.7975956305765248 ind=0.006978706827625781
X6 nt_p_1 nt_c_1 rl_admittance res=1.555726829308897 ind=0.0005181830411010667
* Transfer network from port 2 to port 1
R1_2 nt_p_2 nt_c_1 3.426694989774083
X7 nt_n_2 nt_c_1 rl_admittance res=5.0675924306232725 ind=4.37270294104299e-07
X8 nt_n_2 nt_c_1 rl_admittance res=8.513155152907448 ind=3.254123336075868e-06
X9 nt_p_2 nt_c_1 rl_admittance res=29.19841415943021 ind=2.4511341867419552e-05
X10 nt_n_2 nt_c_1 rl_admittance res=6.835930685348445 ind=0.00023235621768863526
X11 nt_n_2 nt_c_1 rl_admittance res=0.9997197099492963 ind=0.0038811569447894326
X12 nt_p_2 nt_c_1 rl_admittance res=0.8808329569905541 ind=0.0002933887182225766
* Transfer network from port 3 to port 1
R1_3 nt_p_3 nt_c_1 4.441547277752228
X13 nt_n_3 nt_c_1 rl_admittance res=9.905803881729998 ind=8.547478582785004e-07
X14 nt_n_3 nt_c_1 rl_admittance res=6.657668273708107 ind=2.544870063354409e-06
X15 nt_p_3 nt_c_1 rl_admittance res=24.950549841456667 ind=2.094536551213744e-05
X16 nt_n_3 nt_c_1 rl_admittance res=5.320492058717085 ind=0.00018084580840698028
X17 nt_n_3 nt_c_1 rl_admittance res=0.7658650925023123 ind=0.0029732760022185686
X18 nt_p_3 nt_c_1 rl_admittance res=0.6758614717322284 ind=0.00022511661185455517
* Transfer network from port 4 to port 1
R1_4 nt_p_4 nt_c_1 255.40275618332888
X19 nt_n_4 nt_c_1 rl_admittance res=1134.2397565357935 ind=9.787080526209458e-05
X20 nt_n_4 nt_c_1 rl_admittance res=147.65379975650816 ind=5.644014079595739e-05
X21 nt_p_4 nt_c_1 rl_admittance res=239.05992722473442 ind=0.00020068485812313897
X22 nt_n_4 nt_c_1 rl_admittance res=91.00100322070332 ind=0.003093163153270935
X23 nt_n_4 nt_c_1 rl_admittance res=16.831908392482656 ind=0.06534559387136306
X24 nt_p_4 nt_c_1 rl_admittance res=14.294722426174646 ind=0.004761300376738599
* Transfer network from port 5 to port 1
R1_5 nt_n_5 nt_c_1 31.895342935666037
X25 nt_p_5 nt_c_1 rl_admittance res=8.70792321243188 ind=7.513856325792605e-07
X26 nt_n_5 nt_c_1 rl_admittance res=10.476397025500848 ind=4.004565572499293e-06
X27 nt_p_5 nt_c_1 rl_admittance res=47.79808687651375 ind=4.0125304122397295e-05
X28 nt_n_5 nt_c_1 rl_admittance res=8.158140232045698 ind=0.00027729868761754427
X29 nt_n_5 nt_c_1 rl_admittance res=1.116984773206068 ind=0.004336408661956513
X30 nt_p_5 nt_c_1 rl_admittance res=0.9911881113390945 ind=0.0003301459228964249
* Transfer network from port 6 to port 1
R1_6 nt_n_6 nt_c_1 21.076833559021495
X31 nt_p_6 nt_c_1 rl_admittance res=6.109993407294386 ind=5.27216553177767e-07
X32 nt_n_6 nt_c_1 rl_admittance res=7.198365463670849 ind=2.7515496447793397e-06
X33 nt_p_6 nt_c_1 rl_admittance res=28.392200304187178 ind=2.383454540456337e-05
X34 nt_n_6 nt_c_1 rl_admittance res=5.830295211371626 ind=0.00019817423635175733
X35 nt_n_6 nt_c_1 rl_admittance res=0.8296557158751231 ind=0.003220926837199494
X36 nt_p_6 nt_c_1 rl_admittance res=0.7329681351740535 ind=0.00024413775616596723
* Transfer network from port 7 to port 1
R1_7 nt_n_7 nt_c_1 20.442005627247223
X37 nt_p_7 nt_c_1 rl_admittance res=20.902369937839318 ind=1.8036149464118827e-06
X38 nt_p_7 nt_c_1 rl_admittance res=418.1033890288166 ind=0.0001598185362176108
X39 nt_n_7 nt_c_1 rl_admittance res=487.0298192931957 ind=0.00040884940994192836
X40 nt_p_7 nt_c_1 rl_admittance res=111.29034794141766 ind=0.003782806687660541
X41 nt_p_7 nt_c_1 rl_admittance res=16.502908991013452 ind=0.06406833755728226
X42 nt_n_7 nt_c_1 rl_admittance res=14.52602462237651 ind=0.004838342742521081
* Transfer network from port 8 to port 1
R1_8 nt_n_8 nt_c_1 21.135208598873287
X43 nt_p_8 nt_c_1 rl_admittance res=27.412261434985673 ind=2.365337738549323e-06
X44 nt_p_8 nt_c_1 rl_admittance res=76.18582272880558 ind=2.9121760283585987e-05
X45 nt_n_8 nt_c_1 rl_admittance res=288.32487675917 ind=0.00024204155693308856
X46 nt_p_8 nt_c_1 rl_admittance res=64.56543883182214 ind=0.002194606974661626
X47 nt_p_8 nt_c_1 rl_admittance res=9.555668361820281 ind=0.0370974466697915
X48 nt_n_8 nt_c_1 rl_admittance res=8.406102610189041 ind=0.002799913026048667
* Transfer network from port 9 to port 1
R1_9 nt_p_9 nt_c_1 6.008260165842241
X49 nt_n_9 nt_c_1 rl_admittance res=206.56807492333104 ind=1.7824259569188454e-05
X50 nt_n_9 nt_c_1 rl_admittance res=4.369492309650421 ind=1.670222923962732e-06
X51 nt_p_9 nt_c_1 rl_admittance res=11.421088765188914 ind=9.58771971974635e-06
X52 nt_n_9 nt_c_1 rl_admittance res=3.9354441554419886 ind=0.00013376743577041337
X53 nt_n_9 nt_c_1 rl_admittance res=0.6931964771770818 ind=0.0026911586264872704
X54 nt_p_9 nt_c_1 rl_admittance res=0.5965167860048198 ind=0.00019868840494132633
* Transfer network from port 10 to port 1
R1_10 nt_n_10 nt_c_1 36.326812927233185
X55 nt_p_10 nt_c_1 rl_admittance res=13.452724127200316 ind=1.160803027500257e-06
X56 nt_n_10 nt_c_1 rl_admittance res=37.86815320119619 ind=1.4474967131783496e-05
X57 nt_n_10 nt_c_1 rl_admittance res=49.36951526516557 ind=4.144447913800248e-05
X58 nt_n_10 nt_c_1 rl_admittance res=106.29908651629562 ind=0.003613151569781383
X59 nt_n_10 nt_c_1 rl_admittance res=6.579332639499831 ind=0.0255425818974497
X60 nt_p_10 nt_c_1 rl_admittance res=6.201359946230818 ind=0.002065555144618637
* Transfer network from port 11 to port 1
R1_11 nt_n_11 nt_c_1 16.220957163938962
X61 nt_p_11 nt_c_1 rl_admittance res=5.28468649405648 ind=4.5600281576331894e-07
X62 nt_n_11 nt_c_1 rl_admittance res=14.496564596447781 ind=5.541260355171731e-06
X63 nt_n_11 nt_c_1 rl_admittance res=15.875665140189273 ind=1.3327225701337477e-05
X64 nt_p_11 nt_c_1 rl_admittance res=18.99926218067671 ind=0.0006457930752046163
X65 nt_p_11 nt_c_1 rl_admittance res=8.102047186888242 ind=0.03145413298693274
X66 nt_n_11 nt_c_1 rl_admittance res=5.825308378502527 ind=0.0019402995140637318
* Transfer network from port 12 to port 1
R1_12 nt_n_12 nt_c_1 34.84890712168378
X67 nt_p_12 nt_c_1 rl_admittance res=37.191884769599184 ind=3.209197782603766e-06
X68 nt_p_12 nt_c_1 rl_admittance res=83.01733110565019 ind=3.173308010924376e-05
X69 nt_n_12 nt_c_1 rl_admittance res=112.42272148507507 ind=9.437607621222066e-05
X70 nt_n_12 nt_c_1 rl_admittance res=41.382723878587186 ind=0.0014066165443559586
X71 nt_n_12 nt_c_1 rl_admittance res=4.487320520567812 ind=0.017420878100704047
X72 nt_p_12 nt_c_1 rl_admittance res=4.070472154262086 ind=0.0013557969174766587
* Transfer network from port 13 to port 1
R1_13 nt_n_13 nt_c_1 16.3478467890042
X73 nt_p_13 nt_c_1 rl_admittance res=9.30808184900769 ind=8.031718697554935e-07
X74 nt_n_13 nt_c_1 rl_admittance res=190.23771085704544 ind=7.271768964414354e-05
X75 nt_n_13 nt_c_1 rl_admittance res=22.239444620974364 ind=1.8669460165534045e-05
X76 nt_p_13 nt_c_1 rl_admittance res=22.22614011959369 ind=0.0007554760411885568
X77 nt_p_13 nt_c_1 rl_admittance res=9.432199066797386 ind=0.03661810860425445
X78 nt_n_13 nt_c_1 rl_admittance res=6.800268485565257 ind=0.0022650401971400893
* Transfer network from port 14 to port 1
R1_14 nt_n_14 nt_c_1 14.555956665707876
X79 nt_p_14 nt_c_1 rl_admittance res=8.98925428764408 ind=7.756610106178191e-07
X80 nt_p_14 nt_c_1 rl_admittance res=91.04055464134191 ind=3.4799928823862905e-05
X81 nt_n_14 nt_c_1 rl_admittance res=19.674947078207946 ind=1.651662831495207e-05
X82 nt_n_14 nt_c_1 rl_admittance res=18.36911827518103 ind=0.0006243742134255845
X83 nt_n_14 nt_c_1 rl_admittance res=1.4270106482155747 ind=0.005540005095919582
X84 nt_p_14 nt_c_1 rl_admittance res=1.3288974800799649 ind=0.0004426304956412455
* Transfer network from port 15 to port 1
R1_15 nt_p_15 nt_c_1 38.75487733078962
X85 nt_n_15 nt_c_1 rl_admittance res=69.80399782301572 ind=6.023218140684573e-06
X86 nt_n_15 nt_c_1 rl_admittance res=73.17510229100023 ind=2.7970923084088108e-05
X87 nt_p_15 nt_c_1 rl_admittance res=297.14260325091504 ind=0.0002494438188282867
X88 nt_n_15 nt_c_1 rl_admittance res=64.73140214301571 ind=0.002200248138833562
X89 nt_n_15 nt_c_1 rl_admittance res=9.381582334077214 ind=0.03642160204170061
X90 nt_p_15 nt_c_1 rl_admittance res=8.273805721497194 ind=0.002755847446655783
* Transfer network from port 16 to port 1
R1_16 nt_n_16 nt_c_1 23.87622256925236
X91 nt_p_16 nt_c_1 rl_admittance res=26.837078504804023 ind=2.315706594670341e-06
X92 nt_p_16 nt_c_1 rl_admittance res=136.55084304699977 ind=5.2196075008490575e-05
X93 nt_n_16 nt_c_1 rl_admittance res=269.147285290839 ind=0.00022594244627223949
X94 nt_p_16 nt_c_1 rl_admittance res=83.20287728414604 ind=0.0028281015060600202
X95 nt_p_16 nt_c_1 rl_admittance res=13.335713205362934 ind=0.05177250723939369
X96 nt_n_16 nt_c_1 rl_admittance res=11.62892373205639 ind=0.003873373493781197

* Port network for port 2
R_ref_2 p2 a2 50.0
H_b_2 a2 0 V_c_2 14.142135623730951
* Differential incident wave a sources for transfer from port 2
H_p_2 nt_p_2 nts_p_2 H_b_2 3.5355339059327378
E_p_2 nts_p_2 0 p2 0 0.07071067811865475
E_n_2 0 nt_n_2 nt_p_2 0 1
* Current sensor on center node for transfer to port 2
V_c_2 nt_c_2 0 0
* Transfer network from port 1 to port 2
R2_1 nt_p_1 nt_c_2 3.4271018314698125
X97 nt_n_1 nt_c_2 rl_admittance res=5.068597789467925 ind=4.373570440873926e-07
X98 nt_n_1 nt_c_2 rl_admittance res=8.51316124170822 ind=3.2541256634983484e-06
X99 nt_p_1 nt_c_2 rl_admittance res=29.201049666010988 ind=2.4513554309589955e-05
X100 nt_n_1 nt_c_2 rl_admittance res=6.834499729406777 ind=0.00023230757888207193
X101 nt_n_1 nt_c_2 rl_admittance res=0.9995213821731511 ind=0.0038803869877524055
X102 nt_p_1 nt_c_2 rl_admittance res=0.8806563905015528 ind=0.0002933299072806402
* Transfer network from port 2 to port 2
R2_2 nt_p_2 nt_c_2 27.215048698946276
X103 nt_n_2 nt_c_2 rl_admittance res=1.1073020043855104 ind=9.55464117820502e-08
X104 nt_n_2 nt_c_2 rl_admittance res=6.025363975621816 ind=2.303173990048268e-06
X105 nt_p_2 nt_c_2 rl_admittance res=18.189006641347113 ind=1.5269218306872734e-05
X106 nt_n_2 nt_c_2 rl_admittance res=3.473720253045889 ind=0.00011807324217551069
X107 nt_n_2 nt_c_2 rl_admittance res=0.4875495635633539 ind=0.0018927869038902307
X108 nt_p_2 nt_c_2 rl_admittance res=0.43153898353159414 ind=0.00014373743425084593
* Transfer network from port 3 to port 2
R2_3 nt_p_3 nt_c_2 2.971640910246832
X109 nt_n_3 nt_c_2 rl_admittance res=10.136476182596157 ind=8.746520132046011e-07
X110 nt_n_3 nt_c_2 rl_admittance res=3.4945263433776206 ind=1.3357702894247505e-06
X111 nt_p_3 nt_c_2 rl_admittance res=12.99674996707837 ind=1.0910448076699532e-05
X112 nt_n_3 nt_c_2 rl_admittance res=2.5738351952249046 ind=8.748576286739586e-05
X113 nt_n_3 nt_c_2 rl_admittance res=0.3552120716128951 ind=0.0013790203242900459
X114 nt_p_3 nt_c_2 rl_admittance res=0.3149503526475093 ind=0.00010490397700683686
* Transfer network from port 4 to port 2
R2_4 nt_p_4 nt_c_2 31.78444946680438
X115 nt_n_4 nt_c_2 rl_admittance res=36.467565811131365 ind=3.1466980515518764e-06
X116 nt_n_4 nt_c_2 rl_admittance res=85.18167976491611 ind=3.256039470095731e-05
X117 nt_p_4 nt_c_2 rl_admittance res=111.0093975468776 ind=9.318962594716824e-05
X118 nt_n_4 nt_c_2 rl_admittance res=33.37824745077181 ind=0.001134540955390238
X119 nt_n_4 nt_c_2 rl_admittance res=5.3067391526186425 ind=0.020602062069393863
X120 nt_p_4 nt_c_2 rl_admittance res=4.606370196687675 ind=0.0015342943709579747
* Transfer network from port 5 to port 2
R2_5 nt_p_5 nt_c_2 6.175188687232657
X121 nt_p_5 nt_c_2 rl_admittance res=358.3751952847086 ind=3.092332881682761e-05
X122 nt_n_5 nt_c_2 rl_admittance res=5.191885744686813 ind=1.9845798950645147e-06
X123 nt_p_5 nt_c_2 rl_admittance res=21.010543110538933 ind=1.7637827937865863e-05
X124 nt_n_5 nt_c_2 rl_admittance res=3.71434145604034 ind=0.0001262520601297817
X125 nt_n_5 nt_c_2 rl_admittance res=0.5012913500972411 ind=0.0019461358873193117
X126 nt_p_5 nt_c_2 rl_admittance res=0.4455615195213491 ind=0.00014840807449836824
* Transfer network from port 6 to port 2
R2_6 nt_n_6 nt_c_2 29.656860802897047
X127 nt_p_6 nt_c_2 rl_admittance res=3.7473182356940384 ind=3.233470271054931e-07
X128 nt_n_6 nt_c_2 rl_admittance res=3.536594751271808 ind=1.3518507890023107e-06
X129 nt_p_6 nt_c_2 rl_admittance res=12.894988529656187 ind=1.0825021883072864e-05
X130 nt_n_6 nt_c_2 rl_admittance res=2.5961925129527197 ind=8.824569769178377e-05
X131 nt_n_6 nt_c_2 rl_admittance res=0.3593573131894268 ind=0.0013951131680866357
X132 nt_p_6 nt_c_2 rl_admittance res=0.3184718481650312 ind=0.0001060769202396176
* Transfer network from port 7 to port 2
R2_7 nt_p_7 nt_c_2 19.57862671120745
X133 nt_n_7 nt_c_2 rl_admittance res=17.339291424840226 ind=1.4961655193662678e-06
X134 nt_p_7 nt_c_2 rl_admittance res=121.93155078285199 ind=4.66079024380154e-05
X135 nt_n_7 nt_c_2 rl_admittance res=389.81518254989777 ind=0.0003272401423042752
X136 nt_p_7 nt_c_2 rl_admittance res=78.92401581686946 ind=0.0026826611684800977
X137 nt_p_7 nt_c_2 rl_admittance res=10.739990381500094 ind=0.041695275026882195
X138 nt_n_7 nt_c_2 rl_admittance res=9.54016463694869 ind=0.003177647534930672
* Transfer network from port 8 to port 2
R2_8 nt_n_8 nt_c_2 12.672289491521822
X139 nt_p_8 nt_c_2 rl_admittance res=16.445137699203475 ind=1.4190111570262898e-06
X140 nt_p_8 nt_c_2 rl_admittance res=46.79986869175787 ind=1.7889083671066902e-05
X141 nt_n_8 nt_c_2 rl_admittance res=186.77727744652282 ind=0.00015679487507642547
X142 nt_p_8 nt_c_2 rl_admittance res=35.85409800256855 ind=0.0012186961781766271
X143 nt_p_8 nt_c_2 rl_admittance res=5.031148035925612 ind=0.0195321498071562
X144 nt_n_8 nt_c_2 rl_admittance res=4.453110666116599 ind=0.00148324653393872
* Transfer network from port 9 to port 2
R2_9 nt_n_9 nt_c_2 260.31799804428647
X145 nt_p_9 nt_c_2 rl_admittance res=6.828857419536567 ind=5.892455901134532e-07
X146 nt_n_9 nt_c_2 rl_admittance res=5.7893005665287705 ind=2.2129395899315316e-06
X147 nt_p_9 nt_c_2 rl_admittance res=24.233856518920355 ind=2.0343719308105136e-05
X148 nt_n_9 nt_c_2 rl_admittance res=7.502140305305653 ind=0.00025500096858010064
X149 nt_n_9 nt_c_2 rl_admittance res=1.4209649297438829 ind=0.00551653413501011
X150 nt_p_9 nt_c_2 rl_admittance res=1.2107795718184295 ind=0.000403287665165892
* Transfer network from port 10 to port 2
R2_10 nt_n_10 nt_c_2 20.197133834987596
X151 nt_p_10 nt_c_2 rl_admittance res=5.807658758110271 ind=5.011288275414735e-07
X152 nt_n_10 nt_c_2 rl_admittance res=12.12620787000606 ind=4.635199911094885e-06
X153 nt_n_10 nt_c_2 rl_admittance res=25.946684239757936 ind=2.178159554330757e-05
X154 nt_n_10 nt_c_2 rl_admittance res=26.887667781773924 ind=0.0009139233669574745
X155 nt_n_10 nt_c_2 rl_admittance res=2.2184932347335518 ind=0.008612734488741045
X156 nt_p_10 nt_c_2 rl_admittance res=2.0564268838409325 ind=0.0006849567137336445
* Transfer network from port 11 to port 2
R2_11 nt_n_11 nt_c_2 7.918338878519459
X157 nt_p_11 nt_c_2 rl_admittance res=2.804584819234166 ind=2.4200084074167417e-07
X158 nt_n_11 nt_c_2 rl_admittance res=8.074230182679806 ind=3.0863458243602065e-06
X159 nt_n_11 nt_c_2 rl_admittance res=8.967694914984396 ind=7.528156653429424e-06
X160 nt_p_11 nt_c_2 rl_admittance res=17.700479963085424 ind=0.0006016469102460426
X161 nt_n_11 nt_c_2 rl_admittance res=15.159194748297127 ind=0.05885170952341521
X162 nt_p_11 nt_c_2 rl_admittance res=68.66293935084344 ind=0.022870320195971617
* Transfer network from port 12 to port 2
R2_12 nt_n_12 nt_c_2 29.11664426525359
X163 nt_p_12 nt_c_2 rl_admittance res=10.20378857427295 ind=8.804602366772522e-07
X164 nt_n_12 nt_c_2 rl_admittance res=24.539650259509724 ind=9.38019419760468e-06
X165 nt_n_12 nt_c_2 rl_admittance res=49.33801805641684 ind=4.141803801529992e-05
X166 nt_n_12 nt_c_2 rl_admittance res=21.861169417307593 ind=0.000743070530387793
X167 nt_n_12 nt_c_2 rl_admittance res=2.328657267447904 ind=0.009040418264883663
X168 nt_p_12 nt_c_2 rl_admittance res=2.116242394603545 ind=0.0007048801236074417
* Transfer network from port 13 to port 2
R2_13 nt_n_13 nt_c_2 11.421720032076328
X169 nt_p_13 nt_c_2 rl_admittance res=4.2383726441497585 ind=3.657189243222225e-07
X170 nt_n_13 nt_c_2 rl_admittance res=11.84971821306551 ind=4.529512721248876e-06
X171 nt_n_13 nt_c_2 rl_admittance res=14.544369084225108 ind=1.2209635801546778e-05
X172 nt_p_13 nt_c_2 rl_admittance res=16.398141295670353 ind=0.0005573798600316797
X173 nt_p_13 nt_c_2 rl_admittance res=4.094280295936041 ind=0.015894999614734652
X174 nt_n_13 nt_c_2 rl_admittance res=3.3281529113701884 ind=0.0011085444850425904
* Transfer network from port 14 to port 2
R2_14 nt_n_14 nt_c_2 7.242411155883905
X175 nt_p_14 nt_c_2 rl_admittance res=4.1470666633677045 ind=3.57840352077781e-07
X176 nt_p_14 nt_c_2 rl_admittance res=450.6412144602605 ind=0.00017225600448170832
X177 nt_n_14 nt_c_2 rl_admittance res=10.087543220682209 ind=8.46824143031942e-06
X178 nt_n_14 nt_c_2 rl_admittance res=8.471116031453525 ind=0.00028793686935545235
X179 nt_n_14 nt_c_2 rl_admittance res=0.6860893656182168 ind=0.002663567077466514
X180 nt_p_14 nt_c_2 rl_admittance res=0.6371702769370905 ind=0.00021222931017339514
* Transfer network from port 15 to port 2
R2_15 nt_p_15 nt_c_2 18.600132053194102
X181 nt_n_15 nt_c_2 rl_admittance res=29.49651970011329 ind=2.5451833431552116e-06
X182 nt_n_15 nt_c_2 rl_admittance res=42.89035011354757 ind=1.639468407307163e-05
X183 nt_p_15 nt_c_2 rl_admittance res=177.24354132907231 ind=0.00014879154092366562
X184 nt_n_15 nt_c_2 rl_admittance res=34.270610499360416 ind=0.0011648727583764146
X185 nt_n_15 nt_c_2 rl_admittance res=4.737238245448991 ind=0.018391119963393498
X186 nt_p_15 nt_c_2 rl_admittance res=4.200171136355528 ind=0.0013989971835534146
* Transfer network from port 16 to port 2
R2_16 nt_p_16 nt_c_2 22.72209443411551
X187 nt_n_16 nt_c_2 rl_admittance res=20.125699156040586 ind=1.7365979031455249e-06
X188 nt_p_16 nt_c_2 rl_admittance res=130.55409438635823 ind=4.990383912101108e-05
X189 nt_n_16 nt_c_2 rl_admittance res=333.52405169379847 ind=0.0002799851391735015
X190 nt_p_16 nt_c_2 rl_admittance res=76.226153452593 ind=0.0025909596689094
X191 nt_p_16 nt_c_2 rl_admittance res=11.124393424129396 ind=0.04318762185534931
X192 nt_n_16 nt_c_2 rl_admittance res=9.8043938061074 ind=0.003265657249645878

* Port network for port 3
R_ref_3 p3 a3 50.0
H_b_3 a3 0 V_c_3 14.142135623730951
* Differential incident wave a sources for transfer from port 3
H_p_3 nt_p_3 nts_p_3 H_b_3 3.5355339059327378
E_p_3 nts_p_3 0 p3 0 0.07071067811865475
E_n_3 0 nt_n_3 nt_p_3 0 1
* Current sensor on center node for transfer to port 3
V_c_3 nt_c_3 0 0
* Transfer network from port 1 to port 3
R3_1 nt_p_1 nt_c_3 4.442087008590788
X193 nt_n_1 nt_c_3 rl_admittance res=9.911001926495722 ind=8.55196384989082e-07
X194 nt_n_1 nt_c_3 rl_admittance res=6.655991374608841 ind=2.5442290746265926e-06
X195 nt_p_1 nt_c_3 rl_admittance res=24.935005968570373 ind=2.0932316817774135e-05
X196 nt_n_1 nt_c_3 rl_admittance res=5.31397025652499 ind=0.00018062412955158804
X197 nt_n_1 nt_c_3 rl_admittance res=0.7646993475848004 ind=0.002968750294725332
X198 nt_p_1 nt_c_3 rl_admittance res=0.6748541871090088 ind=0.0002247811044894568
* Transfer network from port 2 to port 3
R3_2 nt_p_2 nt_c_3 2.971569900092857
X199 nt_n_2 nt_c_3 rl_admittance res=10.136664175582478 ind=8.746682346647014e-07
X200 nt_n_2 nt_c_3 rl_admittance res=3.4944534922571235 ind=1.3357424423425568e-06
X201 nt_p_2 nt_c_3 rl_admittance res=12.995763090869335 ind=1.0909619618687793e-05
X202 nt_n_2 nt_c_3 rl_admittance res=2.572744511403188 ind=8.744869005622014e-05
X203 nt_n_2 nt_c_3 rl_admittance res=0.35502304951783675 ind=0.001378286494187815
X204 nt_p_2 nt_c_3 rl_admittance res=0.3147863868180074 ind=0.00010484936310511116
* Transfer network from port 3 to port 3
R3_3 nt_n_3 nt_c_3 7.468652346684932
X205 nt_n_3 nt_c_3 rl_admittance res=1.7956501549848956 ind=1.5494230882377887e-07
X206 nt_n_3 nt_c_3 rl_admittance res=2.717505872284293 ind=1.0387569727192617e-06
X207 nt_p_3 nt_c_3 rl_admittance res=10.131366838875584 ind=8.505030266916498e-06
X208 nt_n_3 nt_c_3 rl_admittance res=1.9021765117621057 ind=6.465579596886678e-05
X209 nt_n_3 nt_c_3 rl_admittance res=0.26567108394884936 ind=0.0010314002637300298
X210 nt_p_3 nt_c_3 rl_admittance res=0.23524751916744302 ind=7.835647788360088e-05
* Transfer network from port 4 to port 3
R3_4 nt_p_4 nt_c_3 346.660843572243
X211 nt_p_4 nt_c_3 rl_admittance res=172.17319673739743 ind=1.485640871970825e-05
X212 nt_n_4 nt_c_3 rl_admittance res=47.775073283839085 ind=1.826185216447983e-05
X213 nt_p_4 nt_c_3 rl_admittance res=70.71901342956656 ind=5.936685140617127e-05
X214 nt_n_4 nt_c_3 rl_admittance res=23.09065040836576 ind=0.0007848611169153375
X215 nt_n_4 nt_c_3 rl_admittance res=3.797418386310284 ind=0.014742508920872172
X216 nt_p_4 nt_c_3 rl_admittance res=3.2814560527582253 ind=0.0010929906488873298
* Transfer network from port 5 to port 3
R3_5 nt_p_5 nt_c_3 4.394362643272085
X217 nt_p_5 nt_c_3 rl_admittance res=81.97755104507691 ind=7.073644604647527e-06
X218 nt_n_5 nt_c_3 rl_admittance res=3.6065882242888847 ind=1.3786055455910095e-06
X219 nt_p_5 nt_c_3 rl_admittance res=15.46245001522373 ind=1.298034188985665e-05
X220 nt_n_5 nt_c_3 rl_admittance res=2.655540561560113 ind=9.026296333363285e-05
X221 nt_n_5 nt_c_3 rl_admittance res=0.3596076951035335 ind=0.0013960852120456712
X222 nt_p_5 nt_c_3 rl_admittance res=0.31946696626134286 ind=0.00010640837516582115
* Transfer network from port 6 to port 3
R3_6 nt_p_6 nt_c_3 2.6720431580516113
X223 nt_n_6 nt_c_3 rl_admittance res=28.65820112397462 ind=2.47284686081972e-06
X224 nt_n_6 nt_c_3 rl_admittance res=2.4570961128190154 ind=9.392162666006316e-07
X225 nt_p_6 nt_c_3 rl_admittance res=9.460560526501334 ind=7.941905065676146e-06
X226 nt_n_6 nt_c_3 rl_admittance res=1.9352061501719828 ind=6.577848755334868e-05
X227 nt_n_6 nt_c_3 rl_admittance res=0.2705998222849609 ind=0.001050534833981945
X228 nt_p_6 nt_c_3 rl_admittance res=0.23956882495285922 ind=7.979582271665831e-05
* Transfer network from port 7 to port 3
R3_7 nt_p_7 nt_c_3 55.962845556791095
X229 nt_n_7 nt_c_3 rl_admittance res=35.95867998221667 ind=3.1027875241917134e-06
X230 nt_p_7 nt_c_3 rl_admittance res=83.8751714635187 ind=3.2060986540763945e-05
X231 nt_n_7 nt_c_3 rl_admittance res=321.150465819126 ind=0.00026959782184030946
X232 nt_p_7 nt_c_3 rl_admittance res=57.71936809646144 ind=0.001961906092321392
X233 nt_p_7 nt_c_3 rl_admittance res=7.572644209432413 ind=0.029398860872062556
X234 nt_n_7 nt_c_3 rl_admittance res=6.745478485222798 ind=0.002246790689280155
* Transfer network from port 8 to port 3
R3_8 nt_n_8 nt_c_3 10.592435675336304
X235 nt_p_8 nt_c_3 rl_admittance res=13.986457136213804 ind=1.2068575579345043e-06
X236 nt_p_8 nt_c_3 rl_admittance res=37.42749490757148 ind=1.4306527063352484e-05
X237 nt_n_8 nt_c_3 rl_admittance res=152.1325733766379 ind=0.00012771150840055866
X238 nt_p_8 nt_c_3 rl_admittance res=27.73365389838387 ind=0.0009426787981226698
X239 nt_p_8 nt_c_3 rl_admittance res=3.9290282245825114 ind=0.015253450570545935
X240 nt_n_8 nt_c_3 rl_admittance res=3.474526638111167 ind=0.0011572987916669939
* Transfer network from port 9 to port 3
R3_9 nt_n_9 nt_c_3 29.22840445928682
X241 nt_p_9 nt_c_3 rl_admittance res=5.488315862133113 ind=4.735735014264101e-07
X242 nt_n_9 nt_c_3 rl_admittance res=6.331137239882537 ind=2.420054734837593e-06
X243 nt_p_9 nt_c_3 rl_admittance res=60.29259192090297 ind=5.0614130088594865e-05
X244 nt_n_9 nt_c_3 rl_admittance res=13.946876064702046 ind=0.00047406030285123367
X245 nt_n_9 nt_c_3 rl_admittance res=3.474520721891214 ind=0.013488941045552478
X246 nt_p_9 nt_c_3 rl_admittance res=2.833810448856812 ind=0.0009438884054888516
* Transfer network from port 10 to port 3
R3_10 nt_n_10 nt_c_3 10.620604630749224
X247 nt_p_10 nt_c_3 rl_admittance res=4.571422556549285 ind=3.944569957318919e-07
X248 nt_n_10 nt_c_3 rl_admittance res=14.248760434563405 ind=5.446538093979384e-06
X249 nt_n_10 nt_c_3 rl_admittance res=19.371290845052386 ind=1.6261716465958897e-05
X250 nt_n_10 nt_c_3 rl_admittance res=18.3624321332734 ind=0.0006241469485927335
X251 nt_n_10 nt_c_3 rl_admittance res=1.6478226318443407 ind=0.00639725133726555
X252 nt_p_10 nt_c_3 rl_admittance res=1.5185309312186357 ind=0.000505793794335001
* Transfer network from port 11 to port 3
R3_11 nt_n_11 nt_c_3 6.8196966855210635
X253 nt_p_11 nt_c_3 rl_admittance res=2.0087185399670724 ind=1.7332746442596796e-07
X254 nt_n_11 nt_c_3 rl_admittance res=4.804434873621318 ind=1.836478175024025e-06
X255 nt_n_11 nt_c_3 rl_admittance res=6.7600783140684815 ind=5.674917469897799e-06
X256 nt_p_11 nt_c_3 rl_admittance res=19.157960580240328 ind=0.0006511873019124552
X257 nt_n_11 nt_c_3 rl_admittance res=6.260011535323032 ind=0.024302899105603504
X258 nt_p_11 nt_c_3 rl_admittance res=8.89524074043971 ind=0.0029628356414312007
* Transfer network from port 12 to port 3
R3_12 nt_n_12 nt_c_3 14.324588882165326
X259 nt_p_12 nt_c_3 rl_admittance res=7.256362009714163 ind=6.261339272157532e-07
X260 nt_n_12 nt_c_3 rl_admittance res=25.869929638054373 ind=9.888688767651865e-06
X261 nt_n_12 nt_c_3 rl_admittance res=39.40060853628132 ind=3.307583008939711e-05
X262 nt_n_12 nt_c_3 rl_admittance res=14.938444727526132 ind=0.0005077641472401471
X263 nt_n_12 nt_c_3 rl_admittance res=1.7296618924481002 ind=0.006714971405688352
X264 nt_p_12 nt_c_3 rl_admittance res=1.559760413665398 ind=0.0005195265513941417
* Transfer network from port 13 to port 3
R3_13 nt_n_13 nt_c_3 7.516799637098418
X265 nt_p_13 nt_c_3 rl_admittance res=2.791603590195276 ind=2.4088072188496244e-07
X266 nt_n_13 nt_c_3 rl_admittance res=7.3164717063335125 ind=2.7966953367679974e-06
X267 nt_n_13 nt_c_3 rl_admittance res=10.597008870406997 ind=8.895925161426376e-06
X268 nt_p_13 nt_c_3 rl_admittance res=13.23299579714078 ind=0.00044979520618947143
X269 nt_p_13 nt_c_3 rl_admittance res=3.098619128105979 ind=0.012029598925198589
X270 nt_n_13 nt_c_3 rl_admittance res=2.5482235704440046 ind=0.0008487648437127465
* Transfer network from port 14 to port 3
R3_14 nt_n_14 nt_c_3 5.079220420315103
X271 nt_p_14 nt_c_3 rl_admittance res=2.2695209250792634 ind=1.9583147144752005e-07
X272 nt_n_14 nt_c_3 rl_admittance res=11.120576141177501 ind=4.250800752674554e-06
X273 nt_n_14 nt_c_3 rl_admittance res=6.896245020171284 ind=5.7892260301511735e-06
X274 nt_n_14 nt_c_3 rl_admittance res=6.119800324558468 ind=0.00020801463939238384
X275 nt_n_14 nt_c_3 rl_admittance res=0.5273757952991937 ind=0.00204740209687686
X276 nt_p_14 nt_c_3 rl_admittance res=0.4876206831949602 ind=0.0001624171826065321
* Transfer network from port 15 to port 3
R3_15 nt_p_15 nt_c_3 15.403195451324013
X277 nt_n_15 nt_c_3 rl_admittance res=25.62519085376202 ind=2.2111357403944128e-06
X278 nt_n_15 nt_c_3 rl_admittance res=33.23062911411534 ind=1.27022900123926e-05
X279 nt_p_15 nt_c_3 rl_admittance res=140.62851618606658 ind=0.00011805413875298931
X280 nt_n_15 nt_c_3 rl_admittance res=25.50596580441015 ind=0.0008669587237785639
X281 nt_n_15 nt_c_3 rl_admittance res=3.533600816849522 ind=0.013718304454680308
X282 nt_p_15 nt_c_3 rl_admittance res=3.1319661835747667 ind=0.0010431984144359276
* Transfer network from port 16 to port 3
R3_16 nt_p_16 nt_c_3 59.86092277113375
X283 nt_n_16 nt_c_3 rl_admittance res=38.18256802536646 ind=3.294681444627525e-06
X284 nt_p_16 nt_c_3 rl_admittance res=85.30267568638777 ind=3.2606644962412544e-05
X285 nt_n_16 nt_c_3 rl_admittance res=301.85451211906724 ind=0.00025339934903224827
X286 nt_p_16 nt_c_3 rl_admittance res=63.99757853519416 ind=0.0021753051594775104
X287 nt_p_16 nt_c_3 rl_admittance res=8.976440354622612 ind=0.03484874157737536
X288 nt_n_16 nt_c_3 rl_admittance res=7.939415249727489 ind=0.002644468335418227

* Port network for port 4
R_ref_4 p4 a4 50.0
H_b_4 a4 0 V_c_4 14.142135623730951
* Differential incident wave a sources for transfer from port 4
H_p_4 nt_p_4 nts_p_4 H_b_4 3.5355339059327378
E_p_4 nts_p_4 0 p4 0 0.07071067811865475
E_n_4 0 nt_n_4 nt_p_4 0 1
* Current sensor on center node for transfer to port 4
V_c_4 nt_c_4 0 0
* Transfer network from port 1 to port 4
R4_1 nt_p_1 nt_c_4 255.8311912549191
X289 nt_n_1 nt_c_4 rl_admittance res=1115.1400796181651 ind=9.622274033631263e-05
X290 nt_n_1 nt_c_4 rl_admittance res=147.79542892236853 ind=5.649427804183359e-05
X291 nt_p_1 nt_c_4 rl_admittance res=238.47761354923884 ind=0.00020019602028776168
X292 nt_n_1 nt_c_4 rl_admittance res=90.92895745012903 ind=0.0030907142866101033
X293 nt_n_1 nt_c_4 rl_admittance res=16.83832560338357 ind=0.06537050705693537
X294 nt_p_1 nt_c_4 rl_admittance res=14.296862419835863 ind=0.004762013167957735
* Transfer network from port 2 to port 4
R4_2 nt_p_2 nt_c_4 31.77803869277852
X295 nt_n_2 nt_c_4 rl_admittance res=36.42483514484782 ind=3.1430109257088102e-06
X296 nt_n_2 nt_c_4 rl_admittance res=85.18843144068136 ind=3.256297550505058e-05
X297 nt_p_2 nt_c_4 rl_admittance res=110.66776407014355 ind=9.290283314753673e-05
X298 nt_n_2 nt_c_4 rl_admittance res=33.24622056734784 ind=0.0011300533049622777
X299 nt_n_2 nt_c_4 rl_admittance res=5.282849505480601 ind=0.020509316603864253
X300 nt_p_2 nt_c_4 rl_admittance res=4.585961814945389 ind=0.001527496726849807
* Transfer network from port 3 to port 4
R4_3 nt_p_3 nt_c_4 344.6468699589061
X301 nt_p_3 nt_c_4 rl_admittance res=173.59640421194163 ind=1.4979213850445417e-05
X302 nt_n_3 nt_c_4 rl_admittance res=47.77496646534287 ind=1.8261811333488854e-05
X303 nt_p_3 nt_c_4 rl_admittance res=70.53267356008148 ind=5.921042372419033e-05
X304 nt_n_3 nt_c_4 rl_admittance res=22.993152018509367 ind=0.0007815471048019147
X305 nt_n_3 nt_c_4 rl_admittance res=3.778311384976003 ind=0.014668330858576684
X306 nt_p_3 nt_c_4 rl_admittance res=3.265309229520574 ind=0.0010876124489284564
* Transfer network from port 4 to port 4
R4_4 nt_p_4 nt_c_4 1.148347686483825
X307 nt_p_4 nt_c_4 rl_admittance res=45.34175653924879 ind=3.912430505916659e-06
X308 nt_n_4 nt_c_4 rl_admittance res=360.1450323797293 ind=0.00013766416013672966
X309 nt_p_4 nt_c_4 rl_admittance res=498.4730054068423 ind=0.0004184556798356482
X310 nt_p_4 nt_c_4 rl_admittance res=351.2043817543396 ind=0.011937587657964132
X311 nt_p_4 nt_c_4 rl_admittance res=15.615225190474336 ind=0.060622131472764636
X312 nt_n_4 nt_c_4 rl_admittance res=15.002665832661995 ind=0.004997102871360374
* Transfer network from port 5 to port 4
R4_5 nt_p_5 nt_c_4 305.28658479938804
X313 nt_p_5 nt_c_4 rl_admittance res=397.5719565710291 ind=3.4305522544963975e-05
X314 nt_n_5 nt_c_4 rl_admittance res=72.13255236600061 ind=2.7572412076238478e-05
X315 nt_p_5 nt_c_4 rl_admittance res=103.4999829189376 ind=8.688565929457555e-05
X316 nt_n_5 nt_c_4 rl_admittance res=28.48982759315534 ind=0.0009683814665258652
X317 nt_n_5 nt_c_4 rl_admittance res=4.28354930843246 ind=0.016629788310979488
X318 nt_p_5 nt_c_4 rl_admittance res=3.7458208709511776 ind=0.001247661744826751
* Transfer network from port 6 to port 4
R4_6 nt_n_6 nt_c_4 130.17276052528624
X319 nt_p_6 nt_c_4 rl_admittance res=58.97789836327307 ind=5.08906020285258e-06
X320 nt_n_6 nt_c_4 rl_admittance res=42.83089627495795 ind=1.637195805432784e-05
X321 nt_p_6 nt_c_4 rl_admittance res=62.655328599566815 ind=5.25975887160805e-05
X322 nt_n_6 nt_c_4 rl_admittance res=23.213797718387365 ind=0.0007890469468326126
X323 nt_n_6 nt_c_4 rl_admittance res=4.126290241905388 ind=0.016019270070608292
X324 nt_p_6 nt_c_4 rl_admittance res=3.5268345512925405 ind=0.0011747215634642866
* Transfer network from port 7 to port 4
R4_7 nt_p_7 nt_c_4 111.24491078354666
X325 nt_n_7 nt_c_4 rl_admittance res=102.77878857834807 ind=8.868533080473148e-06
X326 nt_p_7 nt_c_4 rl_admittance res=1045.311219755511 ind=0.00039956650296765935
X327 nt_n_7 nt_c_4 rl_admittance res=3619.5689576776654 ind=0.0030385380401107384
X328 nt_p_7 nt_c_4 rl_admittance res=754.9854741563829 ind=0.025662280274554323
X329 nt_p_7 nt_c_4 rl_admittance res=94.05420605709918 ind=0.36514148054926404
X330 nt_n_7 nt_c_4 rl_admittance res=84.04658016386277 ind=0.027994318593066857
* Transfer network from port 8 to port 4
R4_8 nt_n_8 nt_c_4 589.8217544891857
X331 nt_p_8 nt_c_4 rl_admittance res=925.9107891339737 ind=7.989460253992054e-05
X332 nt_p_8 nt_c_4 rl_admittance res=702.7721118496262 ind=0.00026863214496121977
X333 nt_n_8 nt_c_4 rl_admittance res=1054.3688350955952 ind=0.0008851163912624414
X334 nt_p_8 nt_c_4 rl_admittance res=348.5724531940705 ind=0.011848127276687657
X335 nt_p_8 nt_c_4 rl_admittance res=58.606281054849525 ind=0.2275239474230701
X336 nt_n_8 nt_c_4 rl_admittance res=50.484400897904095 ind=0.01681539451052762
* Transfer network from port 9 to port 4
R4_9 nt_n_9 nt_c_4 394.18183777268973
X337 nt_p_9 nt_c_4 rl_admittance res=211.79578882138293 ind=1.8275346357439322e-05
X338 nt_n_9 nt_c_4 rl_admittance res=471.9560468307922 ind=0.0001804035234891358
X339 nt_p_9 nt_c_4 rl_admittance res=5084.275317037917 ind=0.004268122568696082
X340 nt_n_9 nt_c_4 rl_admittance res=176.25421628815994 ind=0.0059909564525234766
X341 nt_n_9 nt_c_4 rl_admittance res=20.949018941621567 ind=0.08132922612471412
X342 nt_p_9 nt_c_4 rl_admittance res=18.78105136886327 ind=0.006255611287308192
* Transfer network from port 10 to port 4
R4_10 nt_p_10 nt_c_4 3870.124715407051
X343 nt_p_10 nt_c_4 rl_admittance res=256.45390472974475 ind=2.2128787166804394e-05
X344 nt_n_10 nt_c_4 rl_admittance res=165.46927781967543 ind=6.325004404186509e-05
X345 nt_p_10 nt_c_4 rl_admittance res=231.0940086453074 ind=0.0001939976677667647
X346 nt_n_10 nt_c_4 rl_admittance res=21.565234088218116 ind=0.000733011561549058
X347 nt_n_10 nt_c_4 rl_admittance res=2.5754852479432873 ind=0.009998664982572758
X348 nt_p_10 nt_c_4 rl_admittance res=2.312947491460691 ind=0.0007703988530972429
* Transfer network from port 11 to port 4
R4_11 nt_p_11 nt_c_4 361.59776710359085
X349 nt_p_11 nt_c_4 rl_admittance res=146.19270922483858 ind=1.2614615289964644e-05
X350 nt_n_11 nt_c_4 rl_admittance res=93.35022353495873 ind=3.568279155928012e-05
X351 nt_p_11 nt_c_4 rl_admittance res=167.29814370774324 ind=0.00014044262718565406
X352 nt_n_11 nt_c_4 rl_admittance res=10.683943750640099 ind=0.0003631518331830959
X353 nt_n_11 nt_c_4 rl_admittance res=1.1973451953665815 ind=0.00464838751708012
X354 nt_p_11 nt_c_4 rl_admittance res=1.0822422275712251 ind=0.00036047431857942245
* Transfer network from port 12 to port 4
R4_12 nt_p_12 nt_c_4 3219.5789624726335
X355 nt_p_12 nt_c_4 rl_admittance res=484.21599527452634 ind=4.178182708305461e-05
X356 nt_n_12 nt_c_4 rl_admittance res=232.3607218052822 ind=8.881906104527706e-05
X357 nt_p_12 nt_c_4 rl_admittance res=314.9536813637502 ind=0.00026439577554303236
X358 nt_n_12 nt_c_4 rl_admittance res=38.85543433040662 ind=0.0013207128880070318
X359 nt_n_12 nt_c_4 rl_admittance res=5.012970601295861 ind=0.019461580550644005
X360 nt_p_12 nt_c_4 rl_admittance res=4.464853201738229 ind=0.0014871577493937862
* Transfer network from port 13 to port 4
R4_13 nt_p_13 nt_c_4 555.8800694949676
X361 nt_p_13 nt_c_4 rl_admittance res=224.17799879419613 ind=1.9343777307756946e-05
X362 nt_n_13 nt_c_4 rl_admittance res=142.73515304539544 ind=5.456000555149655e-05
X363 nt_p_13 nt_c_4 rl_admittance res=277.9833833823242 ind=0.00023336013066810573
X364 nt_n_13 nt_c_4 rl_admittance res=18.124396971549555 ind=0.0006160560312910705
X365 nt_n_13 nt_c_4 rl_admittance res=2.0356091933316787 ind=0.007902733815238231
X366 nt_p_13 nt_c_4 rl_admittance res=1.839667630648829 ind=0.000612758325886996
* Transfer network from port 14 to port 4
R4_14 nt_p_14 nt_c_4 1311.483878639857
X367 nt_p_14 nt_c_4 rl_admittance res=182.92201668145702 ind=1.578389839504408e-05
X368 nt_n_14 nt_c_4 rl_admittance res=87.35004206499298 ind=3.338924349262269e-05
X369 nt_p_14 nt_c_4 rl_admittance res=81.46455245711353 ind=6.83874639372404e-05
X370 nt_n_14 nt_c_4 rl_admittance res=7.177864907707655 ind=0.00024397870865039683
X371 nt_n_14 nt_c_4 rl_admittance res=0.8165416670788398 ind=0.0031700148855259755
X372 nt_p_14 nt_c_4 rl_admittance res=0.7369533970575912 ind=0.0002454651711616404
* Transfer network from port 15 to port 4
R4_15 nt_p_15 nt_c_4 1240.2705636494015
X373 nt_n_15 nt_c_4 rl_admittance res=9490.56182380033 ind=0.0008189176254250962
X374 nt_n_15 nt_c_4 rl_admittance res=683.458499299702 ind=0.00026124958512602496
X375 nt_p_15 nt_c_4 rl_admittance res=1072.1742587674153 ind=0.0009000636012147078
X376 nt_n_15 nt_c_4 rl_admittance res=318.7885345618528 ind=0.010835759100374676
X377 nt_n_15 nt_c_4 rl_admittance res=50.096803862747386 ind=0.19448807129502066
X378 nt_p_15 nt_c_4 rl_admittance res=43.55210810553751 ind=0.01450637952584211
* Transfer network from port 16 to port 4
R4_16 nt_p_16 nt_c_4 168.80055125755732
X379 nt_n_16 nt_c_4 rl_admittance res=159.73395089489873 ind=1.378305628214529e-05
X380 nt_p_16 nt_c_4 rl_admittance res=1900.1215057821237 ind=0.0007263147002828327
X381 nt_n_16 nt_c_4 rl_admittance res=4301.060041847797 ind=0.0036106328413038203
X382 nt_p_16 nt_c_4 rl_admittance res=1013.677217722976 ind=0.03445532365798764
X383 nt_p_16 nt_c_4 rl_admittance res=136.0525788918249 ind=0.5281894576723907
X384 nt_n_16 nt_c_4 rl_admittance res=120.53964366166844 ind=0.040149464513374554

* Port network for port 5
R_ref_5 p5 a5 50.0
H_b_5 a5 0 V_c_5 14.142135623730951
* Differential incident wave a sources for transfer from port 5
H_p_5 nt_p_5 nts_p_5 H_b_5 3.5355339059327378
E_p_5 nts_p_5 0 p5 0 0.07071067811865475
E_n_5 0 nt_n_5 nt_p_5 0 1
* Current sensor on center node for transfer to port 5
V_c_5 nt_c_5 0 0
* Transfer network from port 1 to port 5
R5_1 nt_n_1 nt_c_5 31.88027818598337
X385 nt_p_1 nt_c_5 rl_admittance res=8.706405231904633 ind=7.512546497110285e-07
X386 nt_n_1 nt_c_5 rl_admittance res=10.473483452062679 ind=4.00345186939554e-06
X387 nt_p_1 nt_c_5 rl_admittance res=47.73722522501055 ind=4.007421228095463e-05
X388 nt_n_1 nt_c_5 rl_admittance res=8.150746072159558 ind=0.00027704735694975225
X389 nt_n_1 nt_c_5 rl_admittance res=1.1158416056983416 ind=0.004331970605501774
X390 nt_p_1 nt_c_5 rl_admittance res=0.9901840176824493 ind=0.0003298114783816499
* Transfer network from port 2 to port 5
R5_2 nt_p_2 nt_c_5 6.176106969741236
X391 nt_p_2 nt_c_5 rl_admittance res=355.5644074934104 ind=3.068079273662935e-05
X392 nt_n_2 nt_c_5 rl_admittance res=5.191717692046127 ind=1.984515657539188e-06
X393 nt_p_2 nt_c_5 rl_admittance res=21.003768231588072 ind=1.76321405956298e-05
X394 nt_n_2 nt_c_5 rl_admittance res=3.712331513693361 ind=0.00012618374132682524
X395 nt_n_2 nt_c_5 rl_admittance res=0.5010073491651117 ind=0.0019450333260923084
X396 nt_p_2 nt_c_5 rl_admittance res=0.4453096417631609 ind=0.00014832417880391547
* Transfer network from port 3 to port 5
R5_3 nt_p_3 nt_c_5 4.395897316728365
X397 nt_p_3 nt_c_5 rl_admittance res=81.2991367589738 ind=7.015105876746638e-06
X398 nt_n_3 nt_c_5 rl_admittance res=3.6058935265877383 ind=1.378339999860876e-06
X399 nt_p_3 nt_c_5 rl_admittance res=15.454891170395637 ind=1.2973996427781466e-05
X400 nt_n_3 nt_c_5 rl_admittance res=2.6551686351417776 ind=9.025032139505847e-05
X401 nt_n_3 nt_c_5 rl_admittance res=0.3595421700311713 ind=0.0013958308276546007
X402 nt_p_3 nt_c_5 rl_admittance res=0.3194099276609075 ind=0.00010638937669200368
* Transfer network from port 4 to port 5
R5_4 nt_p_4 nt_c_5 307.1226835927916
X403 nt_p_4 nt_c_5 rl_admittance res=393.04022621256456 ind=3.391449049300327e-05
X404 nt_n_4 nt_c_5 rl_admittance res=72.12796269232923 ind=2.7570657689770624e-05
X405 nt_p_4 nt_c_5 rl_admittance res=103.7220978856346 ind=8.707211928013686e-05
X406 nt_n_4 nt_c_5 rl_admittance res=28.61646379573115 ind=0.0009726858853983434
X407 nt_n_4 nt_c_5 rl_admittance res=4.306912862330906 ind=0.016720491353607824
X408 nt_p_4 nt_c_5 rl_admittance res=3.7657304436927963 ind=0.0012542932451363896
* Transfer network from port 5 to port 5
R5_5 nt_n_5 nt_c_5 4.249427651703761
X409 nt_n_5 nt_c_5 rl_admittance res=1.5963620632442612 ind=1.3774622139569147e-07
X410 nt_n_5 nt_c_5 rl_admittance res=6.399188575275994 ind=2.44606711621412e-06
X411 nt_p_5 nt_c_5 rl_admittance res=25.755835991551702 ind=2.1621383189614715e-05
X412 nt_n_5 nt_c_5 rl_admittance res=3.8256258885943737 ind=0.00013003466575088642
X413 nt_n_5 nt_c_5 rl_admittance res=0.5268053437178427 ind=0.0020451874640206786
X414 nt_p_5 nt_c_5 rl_admittance res=0.4673283146045992 ind=0.00015565818027450432
* Transfer network from port 6 to port 5
R5_6 nt_p_6 nt_c_5 2.8374864745649275
X415 nt_n_6 nt_c_5 rl_admittance res=8.835002731112317 ind=7.623510168852736e-07
X416 nt_n_6 nt_c_5 rl_admittance res=3.5524304778708204 ind=1.3579039392790287e-06
X417 nt_p_6 nt_c_5 rl_admittance res=14.327948842385553 ind=1.2027956395747757e-05
X418 nt_n_6 nt_c_5 rl_admittance res=2.6531687259086194 ind=9.018234362194658e-05
X419 nt_n_6 nt_c_5 rl_admittance res=0.3655497003651206 ind=0.0014191535328534639
X420 nt_p_6 nt_c_5 rl_admittance res=0.3241512884153111 ind=0.00010796863385231477
* Transfer network from port 7 to port 5
R5_7 nt_n_7 nt_c_5 72.67295513225066
X421 nt_p_7 nt_c_5 rl_admittance res=101.41328326147374 ind=8.75070692935997e-06
X422 nt_p_7 nt_c_5 rl_admittance res=245.55958583235517 ind=9.386427996455422e-05
X423 nt_n_7 nt_c_5 rl_admittance res=1158.9695639104827 ind=0.0009729260993364291
X424 nt_p_7 nt_c_5 rl_admittance res=143.05422833526316 ind=0.004862474613967482
X425 nt_p_7 nt_c_5 rl_admittance res=18.993111302236557 ind=0.07373591327670509
X426 nt_n_7 nt_c_5 rl_admittance res=16.963273929786364 ind=0.005650144168222626
* Transfer network from port 8 to port 5
R5_8 nt_p_8 nt_c_5 30.33419019106582
X427 nt_n_8 nt_c_5 rl_admittance res=18.703155043530348 ind=1.6138500123138258e-06
X428 nt_p_8 nt_c_5 rl_admittance res=43.511088012751834 ind=1.6631958931465047e-05
X429 nt_n_8 nt_c_5 rl_admittance res=232.5107838306881 ind=0.00019518701526791748
X430 nt_p_8 nt_c_5 rl_admittance res=37.56495842513276 ind=0.0012768490581688465
X431 nt_p_8 nt_c_5 rl_admittance res=5.056134323220987 ind=0.019629152698562503
X432 nt_n_8 nt_c_5 rl_admittance res=4.492745083145536 ind=0.0014964480050205333
* Transfer network from port 9 to port 5
R5_9 nt_n_9 nt_c_5 16.037885359939207
X433 nt_p_9 nt_c_5 rl_admittance res=8.09322127370093 ind=6.983444890352234e-07
X434 nt_n_9 nt_c_5 rl_admittance res=23.11494137330117 ind=8.835604283471312e-06
X435 nt_n_9 nt_c_5 rl_admittance res=51.08521160672326 ind=4.2884763508892514e-05
X436 nt_p_9 nt_c_5 rl_admittance res=34.41162214857141 ind=0.0011696658048493593
X437 nt_p_9 nt_c_5 rl_admittance res=4.386582608674612 ind=0.01702978883592631
X438 nt_n_9 nt_c_5 rl_admittance res=3.91545081965563 ind=0.0013041622570153458
* Transfer network from port 10 to port 5
R5_10 nt_n_10 nt_c_5 13.773800425530352
X439 nt_p_10 nt_c_5 rl_admittance res=6.240989572100227 ind=5.385198954049437e-07
X440 nt_n_10 nt_c_5 rl_admittance res=21.587179459079618 ind=8.25162271521123e-06
X441 nt_n_10 nt_c_5 rl_admittance res=25.654145398712245 ind=2.1536016468251752e-05
X442 nt_n_10 nt_c_5 rl_admittance res=21.806526760412364 ind=0.0007412132030295965
X443 nt_n_10 nt_c_5 rl_admittance res=1.9128817100190563 ind=0.007426275644578105
X444 nt_p_10 nt_c_5 rl_admittance res=1.765836671268301 ind=0.0005881666364345446
* Transfer network from port 11 to port 5
R5_11 nt_n_11 nt_c_5 7.321133591311336
X445 nt_p_11 nt_c_5 rl_admittance res=2.8579900844826374 ind=2.466090519113015e-07
X446 nt_n_11 nt_c_5 rl_admittance res=10.030158654888988 ind=3.833992539448839e-06
X447 nt_n_11 nt_c_5 rl_admittance res=8.492739703510615 ind=7.1294435761855896e-06
X448 nt_p_11 nt_c_5 rl_admittance res=23.80427237988792 ind=0.0008091174339838808
X449 nt_n_11 nt_c_5 rl_admittance res=5.35398723869027 ind=0.020785490720004553
X450 nt_p_11 nt_c_5 rl_admittance res=6.715484812350994 ind=0.0022368003668599866
* Transfer network from port 12 to port 5
R5_12 nt_n_12 nt_c_5 22.333040120971745
X451 nt_p_12 nt_c_5 rl_admittance res=8.860080318542419 ind=7.645149012507017e-07
X452 nt_n_12 nt_c_5 rl_admittance res=22.663324086468776 ind=8.662975178790346e-06
X453 nt_n_12 nt_c_5 rl_admittance res=47.07774071070063 ind=3.952059144736225e-05
X454 nt_n_12 nt_c_5 rl_admittance res=21.863923961932297 ind=0.0007431641585417214
X455 nt_n_12 nt_c_5 rl_admittance res=2.4086181960191273 ind=0.009350846187977983
X456 nt_p_12 nt_c_5 rl_admittance res=2.1825018898186137 ind=0.0007269499022379344
* Transfer network from port 13 to port 5
R5_13 nt_n_13 nt_c_5 66.09535822212473
X457 nt_p_13 nt_c_5 rl_admittance res=3.808540615256756 ind=3.286297581624305e-07
X458 nt_n_13 nt_c_5 rl_admittance res=4.891638697867124 ind=1.8698115272743267e-06
X459 nt_n_13 nt_c_5 rl_admittance res=23.672553814102564 ind=1.987251965959776e-05
X460 nt_p_13 nt_c_5 rl_admittance res=589.1980388095287 ind=0.020027094198127537
X461 nt_p_13 nt_c_5 rl_admittance res=10.944993094056619 ind=0.04249114580308183
X462 nt_n_13 nt_c_5 rl_admittance res=10.657834959497889 ind=0.0035499222786555926
* Transfer network from port 14 to port 5
R5_14 nt_n_14 nt_c_5 7.825038476174496
X463 nt_p_14 nt_c_5 rl_admittance res=3.194938934596983 ind=2.756835532262156e-07
X464 nt_n_14 nt_c_5 rl_admittance res=17.151541525879527 ind=6.556115861459109e-06
X465 nt_n_14 nt_c_5 rl_admittance res=8.28947068955566 ind=6.958804298829698e-06
X466 nt_n_14 nt_c_5 rl_admittance res=8.416905405770574 ind=0.00028609422692357073
X467 nt_n_14 nt_c_5 rl_admittance res=0.6894064860033335 ind=0.00267644495182597
X468 nt_p_14 nt_c_5 rl_admittance res=0.6397663520845779 ind=0.00021309401346802784
* Transfer network from port 15 to port 5
R5_15 nt_n_15 nt_c_5 156.62620006469487
X469 nt_p_15 nt_c_5 rl_admittance res=38.34534452408443 ind=3.3087270350024637e-06
X470 nt_n_15 nt_c_5 rl_admittance res=45.10139853037611 ind=1.723984948133252e-05
X471 nt_p_15 nt_c_5 rl_admittance res=224.39288740981112 ind=0.0001883722432967434
X472 nt_n_15 nt_c_5 rl_admittance res=36.42375004069911 ind=0.001238058895423356
X473 nt_n_15 nt_c_5 rl_admittance res=4.9128809411278835 ind=0.019073007957949736
X474 nt_p_15 nt_c_5 rl_admittance res=4.366377383461398 ind=0.0014543573258051072
* Transfer network from port 16 to port 5
R5_16 nt_n_16 nt_c_5 206.72927713077235
X475 nt_p_16 nt_c_5 rl_admittance res=1084.9311988320608 ind=9.361608907799962e-05
X476 nt_p_16 nt_c_5 rl_admittance res=249.79317781091478 ind=9.548255546939444e-05
X477 nt_n_16 nt_c_5 rl_admittance res=1612.757292272936 ind=0.001353869601418354
X478 nt_p_16 nt_c_5 rl_admittance res=189.08489884603696 ind=0.0064270768590544685
X479 nt_p_16 nt_c_5 rl_admittance res=26.346624080275454 ind=0.10228405222310137
X480 nt_n_16 nt_c_5 rl_admittance res=23.412686779768123 ind=0.007798321020970262

* Port network for port 6
R_ref_6 p6 a6 50.0
H_b_6 a6 0 V_c_6 14.142135623730951
* Differential incident wave a sources for transfer from port 6
H_p_6 nt_p_6 nts_p_6 H_b_6 3.5355339059327378
E_p_6 nts_p_6 0 p6 0 0.07071067811865475
E_n_6 0 nt_n_6 nt_p_6 0 1
* Current sensor on center node for transfer to port 6
V_c_6 nt_c_6 0 0
* Transfer network from port 1 to port 6
R6_1 nt_n_1 nt_c_6 21.06691569746533
X481 nt_p_1 nt_c_6 rl_admittance res=6.108864305009943 ind=5.271191256725461e-07
X482 nt_n_1 nt_c_6 rl_admittance res=7.197006056631951 ind=2.7510300162645238e-06
X483 nt_p_1 nt_c_6 rl_admittance res=28.376718923177627 ind=2.3821549170575013e-05
X484 nt_n_1 nt_c_6 rl_admittance res=5.829400630568536 ind=0.0001981438291663439
X485 nt_n_1 nt_c_6 rl_admittance res=0.8295038859623511 ind=0.003220337396264683
X486 nt_p_1 nt_c_6 rl_admittance res=0.7328359696977745 ind=0.00024409373435755162
* Transfer network from port 2 to port 6
R6_2 nt_n_2 nt_c_6 29.69716373548692
X487 nt_p_2 nt_c_6 rl_admittance res=3.7478860282998365 ind=3.233960205561556e-07
X488 nt_n_2 nt_c_6 rl_admittance res=3.536224591688803 ind=1.3517092968157486e-06
X489 nt_p_2 nt_c_6 rl_admittance res=12.88792613536277 ind=1.081909317886368e-05
X490 nt_n_2 nt_c_6 rl_admittance res=2.593893117129783 ind=8.816754024095829e-05
X491 nt_n_2 nt_c_6 rl_admittance res=0.35897813869120015 ind=0.0013936411197490528
X492 nt_p_2 nt_c_6 rl_admittance res=0.31814129254793555 ind=0.00010596681844559265
* Transfer network from port 3 to port 6
R6_3 nt_p_3 nt_c_6 2.6731153159930643
X493 nt_n_3 nt_c_6 rl_admittance res=28.850483811302272 ind=2.489438468844635e-06
X494 nt_n_3 nt_c_6 rl_admittance res=2.456211148963489 ind=9.388779923084181e-07
X495 nt_p_3 nt_c_6 rl_admittance res=9.453719734572106 ind=7.936162391135481e-06
X496 nt_n_3 nt_c_6 rl_admittance res=1.934231875790479 ind=6.574537154900383e-05
X497 nt_n_3 nt_c_6 rl_admittance res=0.27044002398493866 ind=0.001049914457814781
X498 nt_p_3 nt_c_6 rl_admittance res=0.23942934996623935 ind=7.974936624926147e-05
* Transfer network from port 4 to port 6
R6_4 nt_n_4 nt_c_6 129.7171789387956
X499 nt_p_4 nt_c_6 rl_admittance res=58.828352316221796 ind=5.0761562361521236e-06
X500 nt_n_4 nt_c_6 rl_admittance res=42.834342813420896 ind=1.6373275481420323e-05
X501 nt_p_4 nt_c_6 rl_admittance res=62.771198327165656 ind=5.2694858468120884e-05
X502 nt_n_4 nt_c_6 rl_admittance res=23.316566794417867 ind=0.00079254011183105
X503 nt_n_4 nt_c_6 rl_admittance res=4.152017321721653 ind=0.016119148900148535
X504 nt_p_4 nt_c_6 rl_admittance res=3.5478571312625253 ind=0.0011817237853295971
* Transfer network from port 5 to port 6
R6_5 nt_p_5 nt_c_6 2.8376298564156617
X505 nt_n_5 nt_c_6 rl_admittance res=8.835333079309075 ind=7.623795218321752e-07
X506 nt_n_5 nt_c_6 rl_admittance res=3.5528301855862914 ind=1.3580567261343321e-06
X507 nt_p_5 nt_c_6 rl_admittance res=14.33257151517205 ind=1.2031837014482473e-05
X508 nt_n_5 nt_c_6 rl_admittance res=2.65386691311443 ind=9.020607530470463e-05
X509 nt_n_5 nt_c_6 rl_admittance res=0.36566086189798375 ind=0.0014195850891696711
X510 nt_p_5 nt_c_6 rl_admittance res=0.32424865483625703 ind=0.00010800106475673601
* Transfer network from port 6 to port 6
R6_6 nt_p_6 nt_c_6 7.602336442369004
X511 nt_n_6 nt_c_6 rl_admittance res=1.2287595445230213 ind=1.0602668915719461e-07
X512 nt_n_6 nt_c_6 rl_admittance res=2.584473628057371 ind=9.87905869618959e-07
X513 nt_p_6 nt_c_6 rl_admittance res=9.212341464436886 ind=7.733531341848174e-06
X514 nt_n_6 nt_c_6 rl_admittance res=1.955573860935685 ind=6.647079478317086e-05
X515 nt_n_6 nt_c_6 rl_admittance res=0.27989181164355514 ind=0.0010866086141336304
X516 nt_p_6 nt_c_6 rl_admittance res=0.24716781382190522 ind=8.232690149428964e-05
* Transfer network from port 7 to port 6
R6_7 nt_n_7 nt_c_6 17.188258397810806
X517 nt_p_7 nt_c_6 rl_admittance res=19.622187959260724 ind=1.6931511397929207e-06
X518 nt_p_7 nt_c_6 rl_admittance res=118.30445869100072 ind=4.522145936183601e-05
X519 nt_n_7 nt_c_6 rl_admittance res=459.10250098449666 ind=0.00038540512140053563
X520 nt_p_7 nt_c_6 rl_admittance res=75.8300841710427 ind=0.0025774971040532454
X521 nt_p_7 nt_c_6 rl_admittance res=9.969290248986363 ind=0.03870322821427358
X522 nt_n_7 nt_c_6 rl_admittance res=8.88466443091033 ind=0.0029593128737239707
* Transfer network from port 8 to port 6
R6_8 nt_p_8 nt_c_6 21.182435195956145
X523 nt_n_8 nt_c_6 rl_admittance res=13.444225668912267 ind=1.1600697160893804e-06
X524 nt_p_8 nt_c_6 rl_admittance res=31.672512952439526 ind=1.2106705640798645e-05
X525 nt_n_8 nt_c_6 rl_admittance res=143.07537549930333 ind=0.0001201082162381823
X526 nt_p_8 nt_c_6 rl_admittance res=28.398929300922067 ind=0.0009652917945631363
X527 nt_p_8 nt_c_6 rl_admittance res=4.018285248301624 ind=0.01559996821347231
X528 nt_n_8 nt_c_6 rl_admittance res=3.55257060725225 ind=0.0011832937546047285
* Transfer network from port 9 to port 6
R6_9 nt_n_9 nt_c_6 12.584347661419756
X529 nt_p_9 nt_c_6 rl_admittance res=6.169783894280551 ind=5.323757296875211e-07
X530 nt_n_9 nt_c_6 rl_admittance res=16.941667069645266 ind=6.47589209560364e-06
X531 nt_n_9 nt_c_6 rl_admittance res=37.08868634588225 ind=3.113502895991376e-05
X532 nt_p_9 nt_c_6 rl_admittance res=17.108904786993605 ind=0.0005815390161315227
X533 nt_p_9 nt_c_6 rl_admittance res=1.9167773090659488 ind=0.007441399314887384
X534 nt_n_9 nt_c_6 rl_admittance res=1.7337451676638136 ind=0.0005774775664654509
* Transfer network from port 10 to port 6
R6_10 nt_n_10 nt_c_6 9.143993409428484
X535 nt_p_10 nt_c_6 rl_admittance res=4.973945784812368 ind=4.291897515357683e-07
X536 nt_n_10 nt_c_6 rl_admittance res=23.347270217430445 ind=8.924411159388098e-06
X537 nt_n_10 nt_c_6 rl_admittance res=21.94253423223518 ind=1.8420211285007973e-05
X538 nt_n_10 nt_c_6 rl_admittance res=16.4022909153053 ind=0.0005575209073839135
X539 nt_n_10 nt_c_6 rl_admittance res=1.6474638317370416 ind=0.006395858387307301
X540 nt_p_10 nt_c_6 rl_admittance res=1.5044841549212906 ind=0.0005011150801016943
* Transfer network from port 11 to port 6
R6_11 nt_n_11 nt_c_6 5.015046140052124
X541 nt_p_11 nt_c_6 rl_admittance res=2.016041184055769 ind=1.739593176734659e-07
X542 nt_n_11 nt_c_6 rl_admittance res=6.209896974194084 ind=2.3737110736728966e-06
X543 nt_n_11 nt_c_6 rl_admittance res=7.155045038403517 ind=6.006482203296314e-06
X544 nt_p_11 nt_c_6 rl_admittance res=21.26491087797425 ind=0.0007228034467467914
X545 nt_n_11 nt_c_6 rl_admittance res=8.932112999248963 ind=0.03467665191920375
X546 nt_p_11 nt_c_6 rl_admittance res=14.471059412242397 ind=0.0048200348756093124
* Transfer network from port 12 to port 6
R6_12 nt_n_12 nt_c_6 14.482093024310377
X547 nt_p_12 nt_c_6 rl_admittance res=6.913390490508408 ind=5.96539744351672e-07
X548 nt_n_12 nt_c_6 rl_admittance res=20.277355109452383 ind=7.750947007353761e-06
X549 nt_n_12 nt_c_6 rl_admittance res=44.237848296959704 ind=3.713657245784417e-05
X550 nt_n_12 nt_c_6 rl_admittance res=17.07271279415689 ind=0.000580308834762923
X551 nt_n_12 nt_c_6 rl_admittance res=2.167939886232808 ind=0.008416473999262477
X552 nt_p_12 nt_c_6 rl_admittance res=1.9373633265019803 ind=0.0006452989055221494
* Transfer network from port 13 to port 6
R6_13 nt_n_13 nt_c_6 7.609477250483986
X553 nt_p_13 nt_c_6 rl_admittance res=2.5878091433936743 ind=2.2329579197796137e-07
X554 nt_n_13 nt_c_6 rl_admittance res=5.481280292444854 ind=2.0951999336140226e-06
X555 nt_n_13 nt_c_6 rl_admittance res=13.143745626259854 ind=1.1033847273503526e-05
X556 nt_p_13 nt_c_6 rl_admittance res=18.962410272436436 ind=0.000644540463028242
X557 nt_p_13 nt_c_6 rl_admittance res=3.083561173162608 ind=0.011971140253411717
X558 nt_n_13 nt_c_6 rl_admittance res=2.677179915779517 ind=0.0008917177515988437
* Transfer network from port 14 to port 6
R6_14 nt_n_14 nt_c_6 5.416791258535574
X559 nt_p_14 nt_c_6 rl_admittance res=1.911173004378084 ind=1.649104960885375e-07
X560 nt_n_14 nt_c_6 rl_admittance res=5.106787718296502 ind=1.9520514765690364e-06
X561 nt_n_14 nt_c_6 rl_admittance res=7.46695038750477 ind=6.268318979785372e-06
X562 nt_n_14 nt_c_6 rl_admittance res=6.20445424783542 ind=0.0002108920625744672
X563 nt_n_14 nt_c_6 rl_admittance res=0.571529611556754 ind=0.002218818033665461
X564 nt_p_14 nt_c_6 rl_admittance res=0.5257680902261669 ind=0.00017512335891791713
* Transfer network from port 15 to port 6
R6_15 nt_n_15 nt_c_6 32.49583517629983
X565 nt_p_15 nt_c_6 rl_admittance res=17.278689423233786 ind=1.4909363192227e-06
X566 nt_n_15 nt_c_6 rl_admittance res=31.592043058687516 ind=1.2075946309574601e-05
X567 nt_p_15 nt_c_6 rl_admittance res=135.98426822980082 ind=0.00011415540820031207
X568 nt_n_15 nt_c_6 rl_admittance res=26.015429164729447 ind=0.0008842756020360416
X569 nt_n_15 nt_c_6 rl_admittance res=3.6255014799800502 ind=0.014075085353756404
X570 nt_p_15 nt_c_6 rl_admittance res=3.2106768932470877 ind=0.0010694154559735766
* Transfer network from port 16 to port 6
R6_16 nt_n_16 nt_c_6 22.955111404830877
X571 nt_p_16 nt_c_6 rl_admittance res=28.40240594516574 ind=2.450774913519399e-06
X572 nt_p_16 nt_c_6 rl_admittance res=104.25697461080962 ind=3.985185843979804e-05
X573 nt_n_16 nt_c_6 rl_admittance res=512.6736198313398 ind=0.00043037674215724186
X574 nt_p_16 nt_c_6 rl_admittance res=103.35277834218972 ind=0.003513005290512102
X575 nt_p_16 nt_c_6 rl_admittance res=14.418064649277627 ind=0.05597446082843059
X576 nt_n_16 nt_c_6 rl_admittance res=12.768267125299547 ind=0.004252867125469362

* Port network for port 7
R_ref_7 p7 a7 50.0
H_b_7 a7 0 V_c_7 14.142135623730951
* Differential incident wave a sources for transfer from port 7
H_p_7 nt_p_7 nts_p_7 H_b_7 3.5355339059327378
E_p_7 nts_p_7 0 p7 0 0.07071067811865475
E_n_7 0 nt_n_7 nt_p_7 0 1
* Current sensor on center node for transfer to port 7
V_c_7 nt_c_7 0 0
* Transfer network from port 1 to port 7
R7_1 nt_n_1 nt_c_7 20.43584806414111
X577 nt_p_1 nt_c_7 rl_admittance res=20.89814451789856 ind=1.8032503451450084e-06
X578 nt_p_1 nt_c_7 rl_admittance res=415.3151555136025 ind=0.00015875274385445998
X579 nt_n_1 nt_c_7 rl_admittance res=482.7615173338529 ind=0.00040526627669545923
X580 nt_p_1 nt_c_7 rl_admittance res=109.67669736344492 ind=0.003727958012004358
X581 nt_p_1 nt_c_7 rl_admittance res=16.194423700875298 ind=0.06287072205138632
X582 nt_n_1 nt_c_7 rl_admittance res=14.261008054620842 ind=0.00475007076029731
* Transfer network from port 2 to port 7
R7_2 nt_p_2 nt_c_7 19.585645761976153
X583 nt_n_2 nt_c_7 rl_admittance res=17.34351026355801 ind=1.4965295527553294e-06
X584 nt_p_2 nt_c_7 rl_admittance res=121.64068869529916 ind=4.649672143758901e-05
X585 nt_n_2 nt_c_7 rl_admittance res=386.4535544603923 ind=0.0003244181392022205
X586 nt_p_2 nt_c_7 rl_admittance res=78.06989162580979 ind=0.0026536291206718373
X587 nt_p_2 nt_c_7 rl_admittance res=10.6039403782163 ind=0.04116709556835146
X588 nt_n_2 nt_c_7 rl_admittance res=9.420964165330178 ind=0.003137944123174636
* Transfer network from port 3 to port 7
R7_3 nt_p_3 nt_c_7 55.9746931597258
X589 nt_n_3 nt_c_7 rl_admittance res=35.95938741979357 ind=3.10284856726918e-06
X590 nt_p_3 nt_c_7 rl_admittance res=83.73192290096355 ind=3.200623028624991e-05
X591 nt_n_3 nt_c_7 rl_admittance res=318.85310477793985 ind=0.000267669244433128
X592 nt_p_3 nt_c_7 rl_admittance res=57.36567847341809 ind=0.0019498840302454537
X593 nt_p_3 nt_c_7 rl_admittance res=7.526429689987763 ind=0.029219444780424427
X594 nt_n_3 nt_c_7 rl_admittance res=6.704216984085745 ind=0.002233047267403776
* Transfer network from port 4 to port 7
R7_4 nt_p_4 nt_c_7 111.32308727646465
X595 nt_n_4 nt_c_7 rl_admittance res=102.89450490147624 ind=8.878517962118554e-06
X596 nt_p_4 nt_c_7 rl_admittance res=1047.4031276335343 ind=0.0004003661273279028
X597 nt_n_4 nt_c_7 rl_admittance res=3620.5841199597376 ind=0.0030393902435766843
X598 nt_p_4 nt_c_7 rl_admittance res=770.7516774483415 ind=0.026198180290638654
X599 nt_p_4 nt_c_7 rl_admittance res=96.71538321166965 ind=0.37547282251640396
X600 nt_n_4 nt_c_7 rl_admittance res=86.35767589330709 ind=0.028764100659428173
* Transfer network from port 5 to port 7
R7_5 nt_n_5 nt_c_7 72.29424652878659
X601 nt_p_5 nt_c_7 rl_admittance res=100.65004633885516 ind=8.68484906131046e-06
X602 nt_p_5 nt_c_7 rl_admittance res=244.48266187444034 ind=9.345262960464824e-05
X603 nt_n_5 nt_c_7 rl_admittance res=1113.7271928014584 ind=0.0009349462549828686
X604 nt_p_5 nt_c_7 rl_admittance res=137.1561435819753 ind=0.004661996181993574
X605 nt_p_5 nt_c_7 rl_admittance res=18.041136631083837 ind=0.07004011427480746
X606 nt_n_5 nt_c_7 rl_admittance res=16.125058241997177 ind=0.005370950452453017
* Transfer network from port 6 to port 7
R7_6 nt_n_6 nt_c_7 17.191796477066347
X607 nt_p_6 nt_c_7 rl_admittance res=19.62809856492641 ind=1.6936611516601243e-06
X608 nt_p_6 nt_c_7 rl_admittance res=118.01634115924978 ind=4.51113274581219e-05
X609 nt_n_6 nt_c_7 rl_admittance res=454.5980825911753 ind=0.00038162377428525287
X610 nt_p_6 nt_c_7 rl_admittance res=75.2728767476913 ind=0.0025585573846035646
X611 nt_p_6 nt_c_7 rl_admittance res=9.892890397601956 ind=0.038406625265636596
X612 nt_n_6 nt_c_7 rl_admittance res=8.81667521397533 ind=0.0029366669576609884
* Transfer network from port 7 to port 7
R7_7 nt_n_7 nt_c_7 1.6171201944676856
X613 nt_n_7 nt_c_7 rl_admittance res=2.4431953711300727 ind=2.1081741933948544e-07
X614 nt_p_7 nt_c_7 rl_admittance res=30.630643570624425 ind=1.1708454768165415e-05
X615 nt_n_7 nt_c_7 rl_admittance res=270.3055515094055 ind=0.00022691478193066764
X616 nt_n_7 nt_c_7 rl_admittance res=503.316041268538 ind=0.017107928244771746
X617 nt_p_7 nt_c_7 rl_admittance res=72.51830671771437 ind=0.28153384087636135
X618 nt_n_7 nt_c_7 rl_admittance res=82.87031807717594 ind=0.027602528046212278
* Transfer network from port 8 to port 7
R7_8 nt_p_8 nt_c_7 30.22525350575004
X619 nt_n_8 nt_c_7 rl_admittance res=28.512753153501688 ind=2.4602965072353944e-06
X620 nt_p_8 nt_c_7 rl_admittance res=460.7122096544607 ind=0.00017610560664334192
X621 nt_n_8 nt_c_7 rl_admittance res=15665.892504129288 ind=0.013151126795115358
X622 nt_n_8 nt_c_7 rl_admittance res=397.5091012443509 ind=0.013511504945465687
X623 nt_n_8 nt_c_7 rl_admittance res=49.69756302544311 ind=0.19293812051088977
X624 nt_p_8 nt_c_7 rl_admittance res=44.409380141490914 ind=0.014791920549029693
* Transfer network from port 9 to port 7
R7_9 nt_n_9 nt_c_7 43.34098624433028
X625 nt_p_9 nt_c_7 rl_admittance res=135.7008183803131 ind=1.1709295405205959e-05
X626 nt_p_9 nt_c_7 rl_admittance res=42.18967351947328 ind=1.6126852932341086e-05
X627 nt_n_9 nt_c_7 rl_admittance res=94.77809752690197 ind=7.956385361686576e-05
X628 nt_p_9 nt_c_7 rl_admittance res=30.350832518878033 ind=0.001031637822616141
X629 nt_p_9 nt_c_7 rl_admittance res=4.710719772826248 ind=0.018288168753008552
X630 nt_n_9 nt_c_7 rl_admittance res=4.120693100940929 ind=0.0013725245603936208
* Transfer network from port 10 to port 7
R7_10 nt_p_10 nt_c_7 119.0852525548607
X631 nt_p_10 nt_c_7 rl_admittance res=267.58652778720796 ind=2.3089394284510286e-05
X632 nt_n_10 nt_c_7 rl_admittance res=72.8348068937175 ind=2.7840846376502346e-05
X633 nt_p_10 nt_c_7 rl_admittance res=591.0916600981726 ind=0.0004962067349458269
X634 nt_n_10 nt_c_7 rl_admittance res=1390.851972014079 ind=0.04727565542386684
X635 nt_p_10 nt_c_7 rl_admittance res=153.19783353909102 ind=0.5947515385058225
X636 nt_n_10 nt_c_7 rl_admittance res=169.34915991943916 ind=0.056406986780544816
* Transfer network from port 11 to port 7
R7_11 nt_p_11 nt_c_7 152.5447962102997
X637 nt_n_11 nt_c_7 rl_admittance res=126.24420940636398 ind=1.0893307489074449e-05
X638 nt_n_11 nt_c_7 rl_admittance res=233.9556306811136 ind=8.942870930124535e-05
X639 nt_p_11 nt_c_7 rl_admittance res=158.5205395943553 ind=0.00013307404702834328
X640 nt_n_11 nt_c_7 rl_admittance res=117.17668610605807 ind=0.00398288584804518
X641 nt_n_11 nt_c_7 rl_admittance res=24.205926242920004 ind=0.09397333853459242
X642 nt_p_11 nt_c_7 rl_admittance res=20.33432788195977 ind=0.006772978174645835
* Transfer network from port 12 to port 7
R7_12 nt_p_12 nt_c_7 179.23371881124368
X643 nt_p_12 nt_c_7 rl_admittance res=396.8167250071125 ind=3.4240355439954695e-05
X644 nt_n_12 nt_c_7 rl_admittance res=118.65879611428133 ind=4.535690358401122e-05
X645 nt_p_12 nt_c_7 rl_admittance res=4224.9012363864285 ind=0.0035466994198965823
X646 nt_p_12 nt_c_7 rl_admittance res=493.3830331368872 ind=0.01677030103554805
X647 nt_p_12 nt_c_7 rl_admittance res=53.1557811082255 ind=0.20636377071565362
X648 nt_n_12 nt_c_7 rl_admittance res=48.19727315027331 ind=0.01605359572340994
* Transfer network from port 13 to port 7
R7_13 nt_p_13 nt_c_7 582.6266455687357
X649 nt_n_13 nt_c_7 rl_admittance res=169.45498141219 ind=1.4621860493708534e-05
X650 nt_p_13 nt_c_7 rl_admittance res=509.87206280720756 ind=0.0001948967859968372
X651 nt_p_13 nt_c_7 rl_admittance res=458.5026565071552 ind=0.00038490156689339295
X652 nt_p_13 nt_c_7 rl_admittance res=736.0134767695079 ind=0.025017413941391925
X653 nt_p_13 nt_c_7 rl_admittance res=35.37058194685749 ind=0.13731726842842
X654 nt_n_13 nt_c_7 rl_admittance res=33.79739382685981 ind=0.011257269582650681
* Transfer network from port 14 to port 7
R7_14 nt_p_14 nt_c_7 549.5562487561955
X655 nt_n_14 nt_c_7 rl_admittance res=58.52920874598412 ind=5.050343861000014e-06
X656 nt_p_14 nt_c_7 rl_admittance res=109.02266659904163 ind=4.1673527284416615e-05
X657 nt_p_14 nt_c_7 rl_admittance res=165.05570538245033 ind=0.00013856015603130523
X658 nt_p_14 nt_c_7 rl_admittance res=1235.6949511703472 ind=0.04200180169852752
X659 nt_p_14 nt_c_7 rl_admittance res=31.726800981946667 ind=0.12317121763387034
X660 nt_n_14 nt_c_7 rl_admittance res=30.96589669454469 ind=0.010314151698938545
* Transfer network from port 15 to port 7
R7_15 nt_n_15 nt_c_7 89.03827137505998
X661 nt_p_15 nt_c_7 rl_admittance res=87.22699561305569 ind=7.526606479847498e-06
X662 nt_n_15 nt_c_7 rl_admittance res=4638.042839613615 ind=0.0017728754107050081
X663 nt_n_15 nt_c_7 rl_admittance res=8000.107418601201 ind=0.006715891035817817
X664 nt_p_15 nt_c_7 rl_admittance res=607.3366990513107 ind=0.020643635044095002
X665 nt_p_15 nt_c_7 rl_admittance res=77.35579159968752 ind=0.3003141428531386
X666 nt_n_15 nt_c_7 rl_admittance res=69.12558658894655 ind=0.023024419198624788
* Transfer network from port 16 to port 7
R7_16 nt_p_16 nt_c_7 6.098861390642815
X667 nt_n_16 nt_c_7 rl_admittance res=5.93016843633702 ind=5.11699891367584e-07
X668 nt_p_16 nt_c_7 rl_admittance res=218.107931353365 ind=8.337098249147047e-05
X669 nt_p_16 nt_c_7 rl_admittance res=3938.9107111513 ind=0.00330661749296025
X670 nt_n_16 nt_c_7 rl_admittance res=733.5304498551596 ind=0.02493301479096262
X671 nt_n_16 nt_c_7 rl_admittance res=127.74314676051668 ind=0.49593020550128053
X672 nt_p_16 nt_c_7 rl_admittance res=110.90214381515392 ind=0.03693939646994019

* Port network for port 8
R_ref_8 p8 a8 50.0
H_b_8 a8 0 V_c_8 14.142135623730951
* Differential incident wave a sources for transfer from port 8
H_p_8 nt_p_8 nts_p_8 H_b_8 3.5355339059327378
E_p_8 nts_p_8 0 p8 0 0.07071067811865475
E_n_8 0 nt_n_8 nt_p_8 0 1
* Current sensor on center node for transfer to port 8
V_c_8 nt_c_8 0 0
* Transfer network from port 1 to port 8
R8_1 nt_n_1 nt_c_8 21.112971246092872
X673 nt_p_1 nt_c_8 rl_admittance res=27.375202802399663 ind=2.3621400387753506e-06
X674 nt_p_1 nt_c_8 rl_admittance res=76.099558207407 ind=2.9088785976514575e-05
X675 nt_n_1 nt_c_8 rl_admittance res=286.36782885719765 ind=0.00024039866393505677
X676 nt_p_1 nt_c_8 rl_admittance res=63.832131806050995 ind=0.002169681554151164
X677 nt_p_1 nt_c_8 rl_admittance res=9.41579237379071 ind=0.03655441380073085
X678 nt_n_1 nt_c_8 rl_admittance res=8.286070109588572 ind=0.002759932481251
* Transfer network from port 2 to port 8
R8_2 nt_n_2 nt_c_8 12.668065459688126
X679 nt_p_2 nt_c_8 rl_admittance res=16.438436995537568 ind=1.418432969513618e-06
X680 nt_p_2 nt_c_8 rl_admittance res=46.7618287547832 ind=1.787454304019753e-05
X681 nt_n_2 nt_c_8 rl_admittance res=186.00934224940687 ind=0.00015615021259421824
X682 nt_p_2 nt_c_8 rl_admittance res=35.69094017638369 ind=0.001213150373644134
X683 nt_p_2 nt_c_8 rl_admittance res=5.003191448465483 ind=0.019423615482491347
X684 nt_n_2 nt_c_8 rl_admittance res=4.428815436743113 ind=0.0014751542547520242
* Transfer network from port 3 to port 8
R8_3 nt_n_3 nt_c_8 10.590598904596666
X685 nt_p_3 nt_c_8 rl_admittance res=13.984795595949285 ind=1.2067141876437638e-06
X686 nt_p_3 nt_c_8 rl_admittance res=37.37859406007089 ind=1.4287834887990074e-05
X687 nt_n_3 nt_c_8 rl_admittance res=151.33185808967005 ind=0.00012703932784889675
X688 nt_p_3 nt_c_8 rl_admittance res=27.60841002646332 ind=0.0009384217051666936
X689 nt_p_3 nt_c_8 rl_admittance res=3.9076250240313657 ind=0.015170358100093378
X690 nt_n_3 nt_c_8 rl_admittance res=3.4559156486309996 ind=0.0011510998247628765
* Transfer network from port 4 to port 8
R8_4 nt_n_4 nt_c_8 594.7340967479709
X691 nt_p_4 nt_c_8 rl_admittance res=923.9791009605651 ind=7.972792183951538e-05
X692 nt_p_4 nt_c_8 rl_admittance res=701.0265144969541 ind=0.000267964896569913
X693 nt_n_4 nt_c_8 rl_admittance res=1052.2042390280224 ind=0.000883299266745766
X694 nt_p_4 nt_c_8 rl_admittance res=350.49167312576157 ind=0.011913362385814228
X695 nt_p_4 nt_c_8 rl_admittance res=59.29733687814808 ind=0.23020679550652784
X696 nt_n_4 nt_c_8 rl_admittance res=51.035184480536664 ind=0.01699885005456029
* Transfer network from port 5 to port 8
R8_5 nt_p_5 nt_c_8 30.315735920223084
X697 nt_n_5 nt_c_8 rl_admittance res=18.690118144061085 ind=1.6127250897903244e-06
X698 nt_p_5 nt_c_8 rl_admittance res=43.44131124024937 ind=1.6605287007878785e-05
X699 nt_n_5 nt_c_8 rl_admittance res=231.08105718976628 ind=0.0001939867953422311
X700 nt_p_5 nt_c_8 rl_admittance res=37.37208468002274 ind=0.001270293196799266
X701 nt_p_5 nt_c_8 rl_admittance res=5.028105680179457 ind=0.01952033863646986
X702 nt_n_5 nt_c_8 rl_admittance res=4.467995071111133 ind=0.001488204246372383
* Transfer network from port 6 to port 8
R8_6 nt_p_6 nt_c_8 21.18073971608277
X703 nt_n_6 nt_c_8 rl_admittance res=13.441685620787654 ind=1.1598505414801956e-06
X704 nt_p_6 nt_c_8 rl_admittance res=31.635871764759692 ind=1.2092699676881759e-05
X705 nt_n_6 nt_c_8 rl_admittance res=142.42394411240792 ind=0.0001195613558045925
X706 nt_p_6 nt_c_8 rl_admittance res=28.299394927474903 ind=0.0009619085784937047
X707 nt_p_6 nt_c_8 rl_admittance res=4.002167926850585 ind=0.015537396821252505
X708 nt_n_6 nt_c_8 rl_admittance res=3.5384866366335954 ind=0.0011786026516498514
* Transfer network from port 7 to port 8
R8_7 nt_p_7 nt_c_8 30.222344639387423
X709 nt_n_7 nt_c_8 rl_admittance res=28.510851805498593 ind=2.4601324445149036e-06
X710 nt_p_7 nt_c_8 rl_admittance res=461.1969888577286 ind=0.0001762909117728578
X711 nt_n_7 nt_c_8 rl_admittance res=16587.099254186363 ind=0.01392445693071558
X712 nt_n_7 nt_c_8 rl_admittance res=391.2364417536999 ind=0.0132982945574171
X713 nt_n_7 nt_c_8 rl_admittance res=48.83728141539594 ind=0.1895982964461241
X714 nt_p_7 nt_c_8 rl_admittance res=43.64822396448839 ind=0.014538393891829055
* Transfer network from port 8 to port 8
R8_8 nt_n_8 nt_c_8 1.3723682551791947
X715 nt_n_8 nt_c_8 rl_admittance res=3.4363381318494763 ind=2.9651330609688143e-07
X716 nt_p_8 nt_c_8 rl_admittance res=41.426188370397185 ind=1.583501344442721e-05
X717 nt_n_8 nt_c_8 rl_admittance res=318.37583631870456 ind=0.00026726858944197074
X718 nt_n_8 nt_c_8 rl_admittance res=292.5391021867265 ind=0.009943529628792918
X719 nt_p_8 nt_c_8 rl_admittance res=376.7543734495892 ind=1.462652820026752
X720 nt_p_8 nt_c_8 rl_admittance res=2269.8124132234866 ind=0.7560313782951168
* Transfer network from port 9 to port 8
R8_9 nt_p_9 nt_c_8 436.8585713920536
X721 nt_n_9 nt_c_8 rl_admittance res=46.54582309643805 ind=4.0163264969205245e-06
X722 nt_p_9 nt_c_8 rl_admittance res=41.91748332487514 ind=1.6022809196712665e-05
X723 nt_n_9 nt_c_8 rl_admittance res=157.75114080895187 ind=0.00013242815590020098
X724 nt_p_9 nt_c_8 rl_admittance res=47.80986246204699 ind=0.0016250777430650398
X725 nt_p_9 nt_c_8 rl_admittance res=8.205872895367728 ind=0.03185720983487573
X726 nt_n_9 nt_c_8 rl_admittance res=7.087059118961634 ind=0.0023605647068245133
* Transfer network from port 10 to port 8
R8_10 nt_p_10 nt_c_8 147.17166302649312
X727 nt_n_10 nt_c_8 rl_admittance res=55.69430434057038 ind=4.805726816499382e-06
X728 nt_p_10 nt_c_8 rl_admittance res=139.75949822606384 ind=5.3422572060179694e-05
X729 nt_p_10 nt_c_8 rl_admittance res=261.648722528202 ind=0.00021964758949043935
X730 nt_p_10 nt_c_8 rl_admittance res=224.74228702421337 ind=0.007639086785880432
X731 nt_p_10 nt_c_8 rl_admittance res=19.593306465670764 ind=0.07606601800867027
X732 nt_n_10 nt_c_8 rl_admittance res=18.081848513477727 ind=0.006022720104149011
* Transfer network from port 11 to port 8
R8_11 nt_p_11 nt_c_8 314.6214406808649
X733 nt_n_11 nt_c_8 rl_admittance res=23.668473768108377 ind=2.042295355687815e-06
X734 nt_p_11 nt_c_8 rl_admittance res=35.24042305946862 ind=1.347052661337179e-05
X735 nt_p_11 nt_c_8 rl_admittance res=90.17759069580005 ind=7.570184264994074e-05
X736 nt_n_11 nt_c_8 rl_admittance res=214.25122086947263 ind=0.007282490944956898
X737 nt_p_11 nt_c_8 rl_admittance res=557.9694733880327 ind=2.1661742537118718
X738 nt_p_11 nt_c_8 rl_admittance res=403.01371443541694 ind=0.13423620922212434
* Transfer network from port 12 to port 8
R8_12 nt_p_12 nt_c_8 215.01422809582698
X739 nt_n_12 nt_c_8 rl_admittance res=136.42605657547463 ind=1.1771874454968835e-05
X740 nt_p_12 nt_c_8 rl_admittance res=1498.8962767805099 ind=0.0005729477808192975
X741 nt_p_12 nt_c_8 rl_admittance res=596.7619325327568 ind=0.000500966787507812
X742 nt_p_12 nt_c_8 rl_admittance res=194.14706793046943 ind=0.006599142158704169
X743 nt_p_12 nt_c_8 rl_admittance res=23.87836279840996 ind=0.09270165695737935
X744 nt_n_12 nt_c_8 rl_admittance res=21.416308081074057 ind=0.0071333652165259595
* Transfer network from port 13 to port 8
R8_13 nt_p_13 nt_c_8 101.30693615271714
X745 nt_n_13 nt_c_8 rl_admittance res=43.198541507281355 ind=3.7274976644959665e-06
X746 nt_p_13 nt_c_8 rl_admittance res=218.96336999047747 ind=8.369797087375762e-05
X747 nt_p_13 nt_c_8 rl_admittance res=104.90729424926907 ind=8.806706212499286e-05
X748 nt_n_13 nt_c_8 rl_admittance res=100.41214041473535 ind=0.003413051745359937
X749 nt_n_13 nt_c_8 rl_admittance res=25.08608500968824 ind=0.09739033059362975
X750 nt_p_13 nt_c_8 rl_admittance res=20.408015664395023 ind=0.006797522174578815
* Transfer network from port 14 to port 8
R8_14 nt_p_14 nt_c_8 70.0097723197763
X751 nt_n_14 nt_c_8 rl_admittance res=47.09741427694446 ind=4.063921965780224e-06
X752 nt_n_14 nt_c_8 rl_admittance res=190.25847801389028 ind=7.272562781612548e-05
X753 nt_p_14 nt_c_8 rl_admittance res=87.0277310592139 ind=7.305761389268089e-05
X754 nt_p_14 nt_c_8 rl_admittance res=73.16112884549693 ind=0.002486778167134688
X755 nt_p_14 nt_c_8 rl_admittance res=6.483674582938194 ind=0.02517121387613892
X756 nt_n_14 nt_c_8 rl_admittance res=5.981300374189886 ind=0.0019922574832842077
* Transfer network from port 15 to port 8
R8_15 nt_n_15 nt_c_8 12.711586780419548
X757 nt_p_15 nt_c_8 rl_admittance res=12.43947642384105 ind=1.0733723338692937e-06
X758 nt_n_15 nt_c_8 rl_admittance res=564.8065450499399 ind=0.0002158952968204381
X759 nt_n_15 nt_c_8 rl_admittance res=4774.502231408228 ind=0.004008075774314187
X760 nt_p_15 nt_c_8 rl_admittance res=287.2914423008192 ind=0.009765159417196245
X761 nt_p_15 nt_c_8 rl_admittance res=39.95545446451792 ind=0.1551168672917799
X762 nt_n_15 nt_c_8 rl_admittance res=35.39879878912849 ind=0.011790667141752595
* Transfer network from port 16 to port 8
R8_16 nt_p_16 nt_c_8 87.8227083694186
X763 nt_n_16 nt_c_8 rl_admittance res=88.2077092990591 ind=7.611229891809238e-06
X764 nt_n_16 nt_c_8 rl_admittance res=5595.777183473928 ind=0.0021389659637536937
X765 nt_p_16 nt_c_8 rl_admittance res=3972.5018464900463 ind=0.0033348164149122096
X766 nt_n_16 nt_c_8 rl_admittance res=450.50755975688014 ind=0.015312945295013591
X767 nt_n_16 nt_c_8 rl_admittance res=59.03413190501685 ind=0.22918496928943424
X768 nt_p_16 nt_c_8 rl_admittance res=52.53108162205311 ind=0.017497104963688347

* Port network for port 9
R_ref_9 p9 a9 50.0
H_b_9 a9 0 V_c_9 14.142135623730951
* Differential incident wave a sources for transfer from port 9
H_p_9 nt_p_9 nts_p_9 H_b_9 3.5355339059327378
E_p_9 nts_p_9 0 p9 0 0.07071067811865475
E_n_9 0 nt_n_9 nt_p_9 0 1
* Current sensor on center node for transfer to port 9
V_c_9 nt_c_9 0 0
* Transfer network from port 1 to port 9
R9_1 nt_p_1 nt_c_9 6.016633088451305
X769 nt_n_1 nt_c_9 rl_admittance res=227.361836157322 ind=1.9618502933231737e-05
X770 nt_n_1 nt_c_9 rl_admittance res=4.364363863302128 ind=1.6682625935517339e-06
X771 nt_p_1 nt_c_9 rl_admittance res=11.399419571942449 ind=9.569528971414776e-06
X772 nt_n_1 nt_c_9 rl_admittance res=3.9061760033856627 ind=0.00013277259872136027
X773 nt_n_1 nt_c_9 rl_admittance res=0.685346871823709 ind=0.002660684534571403
X774 nt_p_1 nt_c_9 rl_admittance res=0.5900691004027991 ind=0.0001965408034020491
* Transfer network from port 2 to port 9
R9_2 nt_n_2 nt_c_9 260.22016190291185
X775 nt_p_2 nt_c_9 rl_admittance res=6.8287563338682435 ind=5.892368676756244e-07
X776 nt_n_2 nt_c_9 rl_admittance res=5.789160317722195 ind=2.2128859803230922e-06
X777 nt_p_2 nt_c_9 rl_admittance res=24.234600659332447 ind=2.0344343995457625e-05
X778 nt_n_2 nt_c_9 rl_admittance res=7.507656641479209 ind=0.0002551884712140191
X779 nt_n_2 nt_c_9 rl_admittance res=1.4228105997679639 ind=0.005523699478416328
X780 nt_p_2 nt_c_9 rl_admittance res=1.2122563107313085 ind=0.0004037795388331526
* Transfer network from port 3 to port 9
R9_3 nt_n_3 nt_c_9 29.182582079994788
X781 nt_p_3 nt_c_9 rl_admittance res=5.487325661097441 ind=4.734880593739921e-07
X782 nt_n_3 nt_c_9 rl_admittance res=6.332512582269192 ind=2.4205804545825204e-06
X783 nt_p_3 nt_c_9 rl_admittance res=60.46651752333416 ind=5.076013630240531e-05
X784 nt_n_3 nt_c_9 rl_admittance res=14.069411912148656 ind=0.00047822534889317063
X785 nt_n_3 nt_c_9 rl_admittance res=3.5417660213393396 ind=0.013750003779797033
X786 nt_p_3 nt_c_9 rl_admittance res=2.8832813371228068 ind=0.0009603662182029463
* Transfer network from port 4 to port 9
R9_4 nt_n_4 nt_c_9 397.36114004551246
X787 nt_p_4 nt_c_9 rl_admittance res=213.36563600630706 ind=1.841080467411499e-05
X788 nt_n_4 nt_c_9 rl_admittance res=462.2143590241299 ind=0.00017667979790736969
X789 nt_p_4 nt_c_9 rl_admittance res=5029.0319402839505 ind=0.004221747129052905
X790 nt_n_4 nt_c_9 rl_admittance res=166.67893372547908 ind=0.0056654884889098195
X791 nt_n_4 nt_c_9 rl_admittance res=19.628699003431645 ind=0.07620342051495008
X792 nt_p_4 nt_c_9 rl_admittance res=17.624303409531002 ind=0.00587032052542005
* Transfer network from port 5 to port 9
R9_5 nt_n_5 nt_c_9 16.043372967839222
X793 nt_p_5 nt_c_9 rl_admittance res=8.095241583531699 ind=6.985188166840974e-07
X794 nt_n_5 nt_c_9 rl_admittance res=23.13053058978661 ind=8.841563206132209e-06
X795 nt_n_5 nt_c_9 rl_admittance res=51.03672729334267 ind=4.284406213470179e-05
X796 nt_p_5 nt_c_9 rl_admittance res=34.40818926805252 ind=0.0011695491197672744
X797 nt_p_5 nt_c_9 rl_admittance res=4.385558687094744 ind=0.017025813721390635
X798 nt_n_5 nt_c_9 rl_admittance res=3.914574875846592 ind=0.0013038704967793906
* Transfer network from port 6 to port 9
R9_6 nt_n_6 nt_c_9 12.585382186416007
X799 nt_p_6 nt_c_9 rl_admittance res=6.170516484425974 ind=5.324389431192903e-07
X800 nt_n_6 nt_c_9 rl_admittance res=16.953617435484347 ind=6.48046008052264e-06
X801 nt_n_6 nt_c_9 rl_admittance res=37.04552979502618 ind=3.109880010974142e-05
X802 nt_p_6 nt_c_9 rl_admittance res=17.088140438994476 ind=0.0005808332270318483
X803 nt_p_6 nt_c_9 rl_admittance res=1.9144400162121713 ind=0.007432325371159792
X804 nt_n_6 nt_c_9 rl_admittance res=1.7316272480726023 ind=0.0005767721276995276
* Transfer network from port 7 to port 9
R9_7 nt_n_7 nt_c_9 43.36283735365662
X805 nt_p_7 nt_c_9 rl_admittance res=135.9643971995141 ind=1.1732038984009809e-05
X806 nt_p_7 nt_c_9 rl_admittance res=42.183507629725206 ind=1.6124496042873372e-05
X807 nt_n_7 nt_c_9 rl_admittance res=94.79320333754501 ind=7.957653456888029e-05
X808 nt_p_7 nt_c_9 rl_admittance res=30.38331946682312 ind=0.0010327420679188248
X809 nt_p_7 nt_c_9 rl_admittance res=4.717939001271842 ind=0.018316195567263376
X810 nt_n_7 nt_c_9 rl_admittance res=4.126773051792862 ind=0.0013745496764762425
* Transfer network from port 8 to port 9
R9_8 nt_p_8 nt_c_9 441.758073145642
X811 nt_n_8 nt_c_9 rl_admittance res=46.61146701841335 ind=4.0219907521780795e-06
X812 nt_p_8 nt_c_9 rl_admittance res=41.92105236147081 ind=1.602417344828152e-05
X813 nt_n_8 nt_c_9 rl_admittance res=157.66515692465433 ind=0.00013235597456968083
X814 nt_p_8 nt_c_9 rl_admittance res=47.78727940164626 ind=0.0016243101351503203
X815 nt_p_8 nt_c_9 rl_admittance res=8.199592910888864 ind=0.03183282939590794
X816 nt_n_8 nt_c_9 rl_admittance res=7.081901264506883 ind=0.0023588467235278526
* Transfer network from port 9 to port 9
R9_9 nt_p_9 nt_c_9 0.9812724990976042
X817 nt_n_9 nt_c_9 rl_admittance res=0.7836113601898872 ind=6.76159289888983e-08
X818 nt_n_9 nt_c_9 rl_admittance res=0.8522224798104779 ind=3.257590175755923e-07
X819 nt_p_9 nt_c_9 rl_admittance res=1.7816914574860987 ind=1.4956856279332603e-06
X820 nt_n_9 nt_c_9 rl_admittance res=0.6004213775462568 ind=2.040858029837338e-05
X821 nt_n_9 nt_c_9 rl_admittance res=0.09889939924944839 ind=0.00038395170807622395
X822 nt_p_9 nt_c_9 rl_admittance res=0.08580764032142775 ind=2.8580894263561867e-05
* Transfer network from port 10 to port 9
R9_10 nt_n_10 nt_c_9 23.825043004743986
X823 nt_p_10 nt_c_9 rl_admittance res=11.074315749074053 ind=9.555759210899873e-07
X824 nt_n_10 nt_c_9 rl_admittance res=122.54471950927072 ind=4.6842284006981605e-05
X825 nt_n_10 nt_c_9 rl_admittance res=22.61891468534344 ind=1.898801583864063e-05
X826 nt_p_10 nt_c_9 rl_admittance res=22.16388408443139 ind=0.0007533599318357211
X827 nt_p_10 nt_c_9 rl_admittance res=5.373789929864104 ind=0.020862369620770396
X828 nt_n_10 nt_c_9 rl_admittance res=4.402140187467334 ind=0.0014662692361668574
* Transfer network from port 11 to port 9
R9_11 nt_n_11 nt_c_9 14.440966670353324
X829 nt_p_11 nt_c_9 rl_admittance res=5.575510187344819 ind=4.810972888563435e-07
X830 nt_n_11 nt_c_9 rl_admittance res=386.35053125638575 ind=0.00014768111905458917
X831 nt_n_11 nt_c_9 rl_admittance res=8.20490846315405 ind=6.887816414724679e-06
X832 nt_p_11 nt_c_9 rl_admittance res=5.79121185693052 ind=0.00019684577636137391
X833 nt_p_11 nt_c_9 rl_admittance res=1.3880610307197438 ind=0.0053887931342703485
X834 nt_n_11 nt_c_9 rl_admittance res=1.1379853768785793 ind=0.00037904130224548633
* Transfer network from port 12 to port 9
R9_12 nt_n_12 nt_c_9 38.52943661273877
X835 nt_p_12 nt_c_9 rl_admittance res=44.71252390816637 ind=3.858135544074277e-06
X836 nt_p_12 nt_c_9 rl_admittance res=83.6332183926051 ind=3.1968500838324206e-05
X837 nt_n_12 nt_c_9 rl_admittance res=170.66015466181736 ind=0.00014326495169298369
X838 nt_n_12 nt_c_9 rl_admittance res=20.866435960342123 ind=0.0007092591132878176
X839 nt_n_12 nt_c_9 rl_admittance res=2.633327191097414 ind=0.010223221582926411
X840 nt_p_12 nt_c_9 rl_admittance res=2.3520365805244605 ind=0.00078341868579752
* Transfer network from port 13 to port 9
R9_13 nt_n_13 nt_c_9 26.46695237615492
X841 nt_p_13 nt_c_9 rl_admittance res=15.26331867892151 ind=1.3170348521731406e-06
X842 nt_p_13 nt_c_9 rl_admittance res=32.56446877021552 ind=1.2447652585760903e-05
X843 nt_n_13 nt_c_9 rl_admittance res=15.65414315152753 ind=1.3141263506076097e-05
X844 nt_p_13 nt_c_9 rl_admittance res=19.558703085878207 ind=0.000664808711660898
X845 nt_n_13 nt_c_9 rl_admittance res=35.59530380462849 ind=0.1381896937594942
X846 nt_n_13 nt_c_9 rl_admittance res=56.833061008871525 ind=0.018930012540660558
* Transfer network from port 14 to port 9
R9_14 nt_n_14 nt_c_9 16.020079821145607
X847 nt_p_14 nt_c_9 rl_admittance res=11.064585468626934 ind=9.547363187243516e-07
X848 nt_p_14 nt_c_9 rl_admittance res=29.32050576134004 ind=1.1207659241466764e-05
X849 nt_n_14 nt_c_9 rl_admittance res=16.468477536373758 ind=1.3824876951394465e-05
X850 nt_n_14 nt_c_9 rl_admittance res=21.001086762068578 ind=0.0007138359518249548
X851 nt_n_14 nt_c_9 rl_admittance res=1.4906857344690223 ind=0.0057872073874850535
X852 nt_p_14 nt_c_9 rl_admittance res=1.3944889939211726 ind=0.00046447778237072775
* Transfer network from port 15 to port 9
R9_15 nt_n_15 nt_c_9 359.09056213214456
X853 nt_p_15 nt_c_9 rl_admittance res=51.33344106108928 ind=4.429438471516436e-06
X854 nt_n_15 nt_c_9 rl_admittance res=50.16418355565128 ind=1.917508108470073e-05
X855 nt_p_15 nt_c_9 rl_admittance res=219.78693731899503 ind=0.00018450566284878428
X856 nt_n_15 nt_c_9 rl_admittance res=61.99520207501404 ind=0.002107243524260316
X857 nt_n_15 nt_c_9 rl_admittance res=10.688016657654574 ind=0.04149350029218196
X858 nt_p_15 nt_c_9 rl_admittance res=9.226619056430529 ind=0.0030732114608231905
* Transfer network from port 16 to port 9
R9_16 nt_n_16 nt_c_9 31.250777969986533
X859 nt_p_16 nt_c_9 rl_admittance res=253.1366790155992 ind=2.1842551783139893e-05
X860 nt_p_16 nt_c_9 rl_admittance res=23.041760505868744 ind=8.80763115668238e-06
X861 nt_n_16 nt_c_9 rl_admittance res=49.9349502995382 ind=4.191914777430742e-05
X862 nt_p_16 nt_c_9 rl_admittance res=16.557708100834045 ind=0.0005628036042185482
X863 nt_p_16 nt_c_9 rl_admittance res=2.624633812143384 ind=0.010189471755084336
X864 nt_n_16 nt_c_9 rl_admittance res=2.28977082972119 ind=0.0007626791475316582

* Port network for port 10
R_ref_10 p10 a10 50.0
H_b_10 a10 0 V_c_10 14.142135623730951
* Differential incident wave a sources for transfer from port 10
H_p_10 nt_p_10 nts_p_10 H_b_10 3.5355339059327378
E_p_10 nts_p_10 0 p10 0 0.07071067811865475
E_n_10 0 nt_n_10 nt_p_10 0 1
* Current sensor on center node for transfer to port 10
V_c_10 nt_c_10 0 0
* Transfer network from port 1 to port 10
R10_1 nt_n_1 nt_c_10 36.202323606178844
X865 nt_p_1 nt_c_10 rl_admittance res=13.434156632723674 ind=1.1592008833101445e-06
X866 nt_n_1 nt_c_10 rl_admittance res=37.90084541186919 ind=1.4487463613258122e-05
X867 nt_n_1 nt_c_10 rl_admittance res=49.26270310226215 ind=4.1354812986059133e-05
X868 nt_n_1 nt_c_10 rl_admittance res=108.86810131095294 ind=0.003700473485164773
X869 nt_n_1 nt_c_10 rl_admittance res=6.673712707178731 ind=0.0259089884526833
X870 nt_p_1 nt_c_10 rl_admittance res=6.293404820681734 ind=0.0020962135430354916
* Transfer network from port 2 to port 10
R10_2 nt_n_2 nt_c_10 20.166513320829775
X871 nt_p_2 nt_c_10 rl_admittance res=5.802005509396096 ind=5.006410223831592e-07
X872 nt_n_2 nt_c_10 rl_admittance res=12.116885370531053 ind=4.631636418764804e-06
X873 nt_n_2 nt_c_10 rl_admittance res=25.92649298429712 ind=2.176464548695759e-05
X874 nt_n_2 nt_c_10 rl_admittance res=26.912942575755434 ind=0.0009147824680517834
X875 nt_n_2 nt_c_10 rl_admittance res=2.2194470711302445 ind=0.008616437515417798
X876 nt_p_2 nt_c_10 rl_admittance res=2.0573908332012034 ind=0.0006852777869462177
* Transfer network from port 3 to port 10
R10_3 nt_n_3 nt_c_10 10.615956202889446
X877 nt_p_3 nt_c_10 rl_admittance res=4.571352201725633 ind=3.944509249843227e-07
X878 nt_n_3 nt_c_10 rl_admittance res=14.26783923724878 ind=5.453830898577413e-06
X879 nt_n_3 nt_c_10 rl_admittance res=19.34483186619832 ind=1.6239504811839132e-05
X880 nt_n_3 nt_c_10 rl_admittance res=18.46353439461803 ind=0.0006275834578446715
X881 nt_n_3 nt_c_10 rl_admittance res=1.6554474719010919 ind=0.0064268528352100784
X882 nt_p_3 nt_c_10 rl_admittance res=1.52566374031015 ind=0.0005081695974882295
* Transfer network from port 4 to port 10
R10_4 nt_p_4 nt_c_10 4281.57610056768
X883 nt_p_4 nt_c_10 rl_admittance res=252.4036607461549 ind=2.1779301409584434e-05
X884 nt_n_4 nt_c_10 rl_admittance res=160.90752825853954 ind=6.150633146602224e-05
X885 nt_p_4 nt_c_10 rl_admittance res=230.45538456604058 ind=0.0001934615587491241
X886 nt_n_4 nt_c_10 rl_admittance res=21.407469775792496 ind=0.0007276490848639106
X887 nt_n_4 nt_c_10 rl_admittance res=2.5558256039141614 ind=0.009922341425883455
X888 nt_p_4 nt_c_10 rl_admittance res=2.2953905699074006 ind=0.0007645509761875811
* Transfer network from port 5 to port 10
R10_5 nt_n_5 nt_c_10 13.780289377306998
X889 nt_p_5 nt_c_10 rl_admittance res=6.244557895852444 ind=5.388277974309951e-07
X890 nt_n_5 nt_c_10 rl_admittance res=21.640927098919516 ind=8.272167559739556e-06
X891 nt_n_5 nt_c_10 rl_admittance res=25.607435851935147 ind=2.1496804966446407e-05
X892 nt_n_5 nt_c_10 rl_admittance res=21.943985503983832 ind=0.0007458854847150961
X893 nt_n_5 nt_c_10 rl_admittance res=1.9218696421550192 ind=0.007461169000067273
X894 nt_p_5 nt_c_10 rl_admittance res=1.7743546157279955 ind=0.00059100380185517
* Transfer network from port 6 to port 10
R10_6 nt_n_6 nt_c_10 9.145220169470765
X895 nt_p_6 nt_c_10 rl_admittance res=4.975920271689777 ind=4.2936012523282654e-07
X896 nt_n_6 nt_c_10 rl_admittance res=23.418702498352808 ind=8.951715895190923e-06
X897 nt_n_6 nt_c_10 rl_admittance res=21.90650376865067 ind=1.8389964607714494e-05
X898 nt_n_6 nt_c_10 rl_admittance res=16.46525626138301 ind=0.0005596611265191705
X899 nt_n_6 nt_c_10 rl_admittance res=1.6524407652922986 ind=0.0064151800632125605
X900 nt_p_6 nt_c_10 rl_admittance res=1.5091429110297137 ind=0.0005026668232242855
* Transfer network from port 7 to port 10
R10_7 nt_p_7 nt_c_10 119.34940159929387
X901 nt_p_7 nt_c_10 rl_admittance res=267.54482773417965 ind=2.3085796087792323e-05
X902 nt_n_7 nt_c_10 rl_admittance res=72.91222426217858 ind=2.7870438890770195e-05
X903 nt_p_7 nt_c_10 rl_admittance res=589.7237117217179 ind=0.0004950583763353496
X904 nt_n_7 nt_c_10 rl_admittance res=1348.599075881446 ind=0.04583946135115457
X905 nt_p_7 nt_c_10 rl_admittance res=156.34266617825523 ind=0.606960549607856
X906 nt_n_7 nt_c_10 rl_admittance res=173.8523113387148 ind=0.05790690093836354
* Transfer network from port 8 to port 10
R10_8 nt_p_8 nt_c_10 147.34782800552475
X907 nt_n_8 nt_c_10 rl_admittance res=55.67555202089754 ind=4.804108724190118e-06
X908 nt_p_8 nt_c_10 rl_admittance res=139.92738421778006 ind=5.348674588452934e-05
X909 nt_p_8 nt_c_10 rl_admittance res=259.7200969687129 ind=0.00021802855634142114
X910 nt_p_8 nt_c_10 rl_admittance res=230.22509205703267 ind=0.007825449681935041
X911 nt_p_8 nt_c_10 rl_admittance res=19.964604178618888 ind=0.07750748673520576
X912 nt_n_8 nt_c_10 rl_admittance res=18.431590811414235 ind=0.006139212616929628
* Transfer network from port 9 to port 10
R10_9 nt_n_9 nt_c_10 23.771784506611073
X913 nt_p_9 nt_c_10 rl_admittance res=11.059565378883827 ind=9.543031473222607e-07
X914 nt_n_9 nt_c_10 rl_admittance res=122.48695907080906 ind=4.682020528442527e-05
X915 nt_n_9 nt_c_10 rl_admittance res=22.60841506621585 ind=1.897920166974403e-05
X916 nt_p_9 nt_c_10 rl_admittance res=22.16350244402422 ind=0.0007533469597144974
X917 nt_p_9 nt_c_10 rl_admittance res=5.38289767656909 ind=0.020897728125782996
X918 nt_n_9 nt_c_10 rl_admittance res=4.408193585610501 ind=0.001468285508046809
* Transfer network from port 10 to port 10
R10_10 nt_p_10 nt_c_10 1.3797436723842311
X919 nt_p_10 nt_c_10 rl_admittance res=3.1039278182042924 ind=2.6783042411675845e-07
X920 nt_n_10 nt_c_10 rl_admittance res=0.5044121501812864 ind=1.9280975377789809e-07
X921 nt_n_10 nt_c_10 rl_admittance res=22.442137715823872 ind=1.8839615973136935e-05
X922 nt_p_10 nt_c_10 rl_admittance res=18.995079973245403 ind=0.0006456509201791988
X923 nt_p_10 nt_c_10 rl_admittance res=0.5363719617778094 ind=0.0020823274201024395
X924 nt_n_10 nt_c_10 rl_admittance res=0.5213875792353918 ind=0.00017366429395611736
* Transfer network from port 11 to port 10
R10_11 nt_n_11 nt_c_10 5.839853704818978
X925 nt_p_11 nt_c_10 rl_admittance res=3.8033698741689417 ind=3.2818358742017774e-07
X926 nt_n_11 nt_c_10 rl_admittance res=194.3611241212275 ind=7.429384972653989e-05
X927 nt_n_11 nt_c_10 rl_admittance res=13.313754656842669 ind=1.1176565622740247e-05
X928 nt_n_11 nt_c_10 rl_admittance res=4.245332514096682 ind=0.00014430067407212295
X929 nt_n_11 nt_c_10 rl_admittance res=0.45786130600559855 ind=0.0017775298114749742
X930 nt_p_11 nt_c_10 rl_admittance res=0.41524995846943985 ind=0.00013831186956669877
* Transfer network from port 12 to port 10
R10_12 nt_n_12 nt_c_10 3.726012727589009
X931 nt_p_12 nt_c_10 rl_admittance res=1.9041204954461164 ind=1.643019521503512e-07
X932 nt_n_12 nt_c_10 rl_admittance res=10.874358367164517 ind=4.156684882614477e-06
X933 nt_n_12 nt_c_10 rl_admittance res=6.405055910408426 ind=5.3768849993948025e-06
X934 nt_n_12 nt_c_10 rl_admittance res=4.241929390509651 ind=0.0001441850004409224
X935 nt_n_12 nt_c_10 rl_admittance res=0.29777198460685905 ind=0.0011560238279980073
X936 nt_p_12 nt_c_10 rl_admittance res=0.2789160601671937 ind=9.29016389937616e-05
* Transfer network from port 13 to port 10
R10_13 nt_n_13 nt_c_10 8.915752658671114
X937 nt_p_13 nt_c_10 rl_admittance res=5.850539196454447 ind=5.048288768534053e-07
X938 nt_p_13 nt_c_10 rl_admittance res=303.6685089888215 ind=0.00011607620955838011
X939 nt_n_13 nt_c_10 rl_admittance res=18.025646762188632 ind=1.5132081754743217e-05
X940 nt_n_13 nt_c_10 rl_admittance res=7.684483910680832 ind=0.00026119890598100135
X941 nt_n_13 nt_c_10 rl_admittance res=0.7615121133586549 ind=0.0029563766702700306
X942 nt_p_13 nt_c_10 rl_admittance res=0.6960254257619903 ind=0.00023183284173689623
* Transfer network from port 14 to port 10
R10_14 nt_n_14 nt_c_10 11.157910956910618
X943 nt_p_14 nt_c_10 rl_admittance res=12.695469893624827 ind=1.0954613912182418e-06
X944 nt_p_14 nt_c_10 rl_admittance res=13.449890823371877 ind=5.141173021034323e-06
X945 nt_n_14 nt_c_10 rl_admittance res=18.273598593049673 ind=1.5340231144627966e-05
X946 nt_n_14 nt_c_10 rl_admittance res=6.2668990488912755 ind=0.00021301458816103526
X947 nt_n_14 nt_c_10 rl_admittance res=0.9823036765194784 ind=0.0038135436343544
X948 nt_p_14 nt_c_10 rl_admittance res=0.8555701225369291 ind=0.0002849741481724942
* Transfer network from port 15 to port 10
R10_15 nt_n_15 nt_c_10 131.25562102584112
X949 nt_p_15 nt_c_10 rl_admittance res=55.40539829365207 ind=4.780797812473511e-06
X950 nt_n_15 nt_c_10 rl_admittance res=167.73071285511378 ind=6.411446955622051e-05
X951 nt_n_15 nt_c_10 rl_admittance res=232.51299104071623 ind=0.00019518886816579327
X952 nt_n_15 nt_c_10 rl_admittance res=245.8359312410426 ind=0.008356068805314464
X953 nt_n_15 nt_c_10 rl_admittance res=19.77497038726349 ind=0.07677128187802326
X954 nt_p_15 nt_c_10 rl_admittance res=18.3591586015201 ind=0.006115086824348621
* Transfer network from port 16 to port 10
R10_16 nt_p_16 nt_c_10 116.50489645067346
X955 nt_p_16 nt_c_10 rl_admittance res=92.0540596318112 ind=7.943122159045854e-06
X956 nt_n_16 nt_c_10 rl_admittance res=46.89829864823165 ind=1.792670817250934e-05
X957 nt_p_16 nt_c_10 rl_admittance res=469.9143225037247 ind=0.00039448137643343886
X958 nt_n_16 nt_c_10 rl_admittance res=360.9488727716896 ind=0.012268807089569138
X959 nt_n_16 nt_c_10 rl_admittance res=227.2349184012618 ind=0.8821816483906747
X960 nt_p_16 nt_c_10 rl_admittance res=144.51121975942291 ind=0.04813394094477874

* Port network for port 11
R_ref_11 p11 a11 50.0
H_b_11 a11 0 V_c_11 14.142135623730951
* Differential incident wave a sources for transfer from port 11
H_p_11 nt_p_11 nts_p_11 H_b_11 3.5355339059327378
E_p_11 nts_p_11 0 p11 0 0.07071067811865475
E_n_11 0 nt_n_11 nt_p_11 0 1
* Current sensor on center node for transfer to port 11
V_c_11 nt_c_11 0 0
* Transfer network from port 1 to port 11
R11_1 nt_n_1 nt_c_11 16.209800578441218
X961 nt_p_1 nt_c_11 rl_admittance res=5.284748893770274 ind=4.5600820008369914e-07
X962 nt_n_1 nt_c_11 rl_admittance res=14.510957543640746 ind=5.546762008142256e-06
X963 nt_n_1 nt_c_11 rl_admittance res=15.86205436590564 ind=1.3315799795131587e-05
X964 nt_p_1 nt_c_11 rl_admittance res=18.797845623774943 ind=0.0006389468399960192
X965 nt_p_1 nt_c_11 rl_admittance res=7.794062345911091 ind=0.030258460347339623
X966 nt_n_1 nt_c_11 rl_admittance res=5.647305726338375 ind=0.0018810102134713836
* Transfer network from port 2 to port 11
R11_2 nt_n_2 nt_c_11 7.921130253253595
X967 nt_p_2 nt_c_11 rl_admittance res=2.805474486304915 ind=2.420776079614155e-07
X968 nt_n_2 nt_c_11 rl_admittance res=8.08351007967573 ind=3.0898930320438936e-06
X969 nt_n_2 nt_c_11 rl_admittance res=8.959838948726286 ind=7.521561765309815e-06
X970 nt_p_2 nt_c_11 rl_admittance res=17.55379539491917 ind=0.0005966610388232306
X971 nt_n_2 nt_c_11 rl_admittance res=16.138948706221544 ind=0.06265535452524892
X972 nt_p_2 nt_c_11 rl_admittance res=98.89911351807642 ind=0.03294141518904213
* Transfer network from port 3 to port 11
R11_3 nt_n_3 nt_c_11 6.80366311392048
X973 nt_p_3 nt_c_11 rl_admittance res=2.0069410647900723 ind=1.7317409039203556e-07
X974 nt_n_3 nt_c_11 rl_admittance res=4.8033373635659595 ind=1.8360586557014506e-06
X975 nt_n_3 nt_c_11 rl_admittance res=6.757706001416716 ind=5.672925972479263e-06
X976 nt_p_3 nt_c_11 rl_admittance res=19.110976170444307 ind=0.0006495902816597579
X977 nt_n_3 nt_c_11 rl_admittance res=6.2942789039737015 ind=0.024435933429619132
X978 nt_p_3 nt_c_11 rl_admittance res=8.974586270097058 ind=0.0029892641294414534
* Transfer network from port 4 to port 11
R11_4 nt_p_4 nt_c_11 363.11116463764375
X979 nt_p_4 nt_c_11 rl_admittance res=145.8969788340487 ind=1.2589097429811798e-05
X980 nt_n_4 nt_c_11 rl_admittance res=92.99510881365889 ind=3.5547050217696406e-05
X981 nt_p_4 nt_c_11 rl_admittance res=168.8414912865917 ind=0.00014173822906042886
X982 nt_n_4 nt_c_11 rl_admittance res=10.670715268968499 ind=0.00036270219141397084
X983 nt_n_4 nt_c_11 rl_admittance res=1.195464246688478 ind=0.004641085213292208
X984 nt_p_4 nt_c_11 rl_admittance res=1.0805764384125707 ind=0.0003599194758680911
* Transfer network from port 5 to port 11
R11_5 nt_n_5 nt_c_11 7.323037134587506
X985 nt_p_5 nt_c_11 rl_admittance res=2.858764798477691 ind=2.466759001081724e-07
X986 nt_n_5 nt_c_11 rl_admittance res=10.047545255591672 ind=3.840638505846187e-06
X987 nt_n_5 nt_c_11 rl_admittance res=8.481970978876786 ind=7.120403499915192e-06
X988 nt_p_5 nt_c_11 rl_admittance res=23.397355051003377 ind=0.0007952861393433098
X989 nt_n_5 nt_c_11 rl_admittance res=5.536640012284952 ind=0.021494593555196236
X990 nt_p_5 nt_c_11 rl_admittance res=7.03959796735211 ind=0.0023447562991967376
* Transfer network from port 6 to port 11
R11_6 nt_n_6 nt_c_11 5.014705520128873
X991 nt_p_6 nt_c_11 rl_admittance res=2.0162450437220176 ind=1.739769082310013e-07
X992 nt_n_6 nt_c_11 rl_admittance res=6.217273703817644 ind=2.376530802384613e-06
X993 nt_n_6 nt_c_11 rl_admittance res=7.14684432952844 ind=5.999597912331242e-06
X994 nt_p_6 nt_c_11 rl_admittance res=20.959987555850596 ind=0.0007124389721675567
X995 nt_n_6 nt_c_11 rl_admittance res=9.421314033893204 ind=0.036575850238604664
X996 nt_p_6 nt_c_11 rl_admittance res=15.96449162319834 ind=0.00531746876321233
* Transfer network from port 7 to port 11
R11_7 nt_p_7 nt_c_11 153.02889834510148
X997 nt_n_7 nt_c_11 rl_admittance res=126.70733581437109 ind=1.0933269546680535e-05
X998 nt_n_7 nt_c_11 rl_admittance res=231.9115790695772 ind=8.864737782898005e-05
X999 nt_p_7 nt_c_11 rl_admittance res=157.60991690861815 ind=0.00013230960195127658
X1000 nt_n_7 nt_c_11 rl_admittance res=115.93925974282442 ind=0.003940825194907572
X1001 nt_n_7 nt_c_11 rl_admittance res=23.745902529493947 ind=0.09218741372750633
X1002 nt_p_7 nt_c_11 rl_admittance res=19.975148675422574 ind=0.006653342406953641
* Transfer network from port 8 to port 11
R11_8 nt_p_8 nt_c_11 315.42782029897904
X1003 nt_n_8 nt_c_11 rl_admittance res=23.674081430561202 ind=2.0427792273178947e-06
X1004 nt_p_8 nt_c_11 rl_admittance res=35.253288977302454 ind=1.347544456479064e-05
X1005 nt_p_8 nt_c_11 rl_admittance res=90.04939477934587 ind=7.559422536918509e-05
X1006 nt_n_8 nt_c_11 rl_admittance res=206.59040864348756 ind=0.007022096649697597
X1007 nt_p_8 nt_c_11 rl_admittance res=3038.7646790862545 ind=11.797229283810571
X1008 nt_p_8 nt_c_11 rl_admittance res=243.318695587868 ind=0.0810448333609291
* Transfer network from port 9 to port 11
R11_9 nt_n_9 nt_c_11 14.452388228348253
X1009 nt_p_9 nt_c_11 rl_admittance res=5.577774388592595 ind=4.812926613057029e-07
X1010 nt_n_9 nt_c_11 rl_admittance res=389.25771529846935 ind=0.00014879237983436957
X1011 nt_n_9 nt_c_11 rl_admittance res=8.204970336839425 ind=6.887868356143364e-06
X1012 nt_p_9 nt_c_11 rl_admittance res=5.793911555177913 ind=0.00019693754026339964
X1013 nt_p_9 nt_c_11 rl_admittance res=1.3894405998036878 ind=0.0053941489595858635
X1014 nt_n_9 nt_c_11 rl_admittance res=1.1390141315174651 ind=0.0003793839608647772
* Transfer network from port 10 to port 11
R11_10 nt_n_10 nt_c_11 5.8425854706386104
X1015 nt_p_10 nt_c_11 rl_admittance res=3.8059775675939815 ind=3.2840859897872583e-07
X1016 nt_n_10 nt_c_11 rl_admittance res=199.51792008223126 ind=7.626501667635792e-05
X1017 nt_n_10 nt_c_11 rl_admittance res=13.302600875583938 ind=1.1167202301018238e-05
X1018 nt_n_10 nt_c_11 rl_admittance res=4.256424740581118 ind=0.0001446777036106455
X1019 nt_n_10 nt_c_11 rl_admittance res=0.458922510852792 ind=0.0017816496687925198
X1020 nt_p_10 nt_c_11 rl_admittance res=0.41622376327827365 ind=0.00013863622544189088
* Transfer network from port 11 to port 11
R11_11 nt_p_11 nt_c_11 1.359445143337768
X1021 nt_p_11 nt_c_11 rl_admittance res=6.818241392417873 ind=5.883295588098387e-07
X1022 nt_n_11 nt_c_11 rl_admittance res=0.5624109956816201 ind=2.1497960657843553e-07
X1023 nt_n_11 nt_c_11 rl_admittance res=15.993108473770384 ind=1.3425816456429096e-05
X1024 nt_n_11 nt_c_11 rl_admittance res=2.6063096652886997 ind=8.858958404153957e-05
X1025 nt_n_11 nt_c_11 rl_admittance res=0.6733758872735448 ind=0.0026142102384657546
X1026 nt_p_11 nt_c_11 rl_admittance res=0.5417777651473749 ind=0.00018045587737901248
* Transfer network from port 12 to port 11
R11_12 nt_n_12 nt_c_11 8.684594823808453
X1027 nt_p_12 nt_c_11 rl_admittance res=6.826278700128559 ind=5.890230786527568e-07
X1028 nt_n_12 nt_c_11 rl_admittance res=101.22496886693561 ind=3.8692885007616814e-05
X1029 nt_n_12 nt_c_11 rl_admittance res=67.89112854537879 ind=5.69929124388165e-05
X1030 nt_n_12 nt_c_11 rl_admittance res=8.767909264375497 ind=0.0002980249987136301
X1031 nt_n_12 nt_c_11 rl_admittance res=1.8858442720703998 ind=0.007321309683599839
X1032 nt_p_12 nt_c_11 rl_admittance res=1.5684290057038517 ind=0.0005224138946602765
* Transfer network from port 13 to port 11
R11_13 nt_n_13 nt_c_11 4.942743431600294
X1033 nt_p_13 nt_c_11 rl_admittance res=2.7187050585181174 ind=2.3459048390259925e-07
X1034 nt_p_13 nt_c_11 rl_admittance res=16.034069062151623 ind=6.128965979150521e-06
X1035 nt_n_13 nt_c_11 rl_admittance res=4.344876941572081 ind=3.6474160379133354e-06
X1036 nt_n_13 nt_c_11 rl_admittance res=21.893974238851477 ind=0.0007441855803505179
X1037 nt_n_13 nt_c_11 rl_admittance res=0.4893396097213679 ind=0.0018997363018149972
X1038 nt_p_13 nt_c_11 rl_admittance res=0.4781190374941207 ind=0.00015925236499718796
* Transfer network from port 14 to port 11
R11_14 nt_n_14 nt_c_11 3.2823218744795186
X1039 nt_p_14 nt_c_11 rl_admittance res=2.6816548240503213 ind=2.3139350878193553e-07
X1040 nt_p_14 nt_c_11 rl_admittance res=5.981349158706653 ind=2.2863494825320597e-06
X1041 nt_n_14 nt_c_11 rl_admittance res=4.5004891096285276 ind=3.7780485794320328e-06
X1042 nt_n_14 nt_c_11 rl_admittance res=3.968894420309045 ind=0.00013490442462868997
X1043 nt_n_14 nt_c_11 rl_admittance res=0.680421259594269 ind=0.0026415621006317938
X1044 nt_p_14 nt_c_11 rl_admittance res=0.5853404793939105 ind=0.00019496578960885713
* Transfer network from port 15 to port 11
R11_15 nt_n_15 nt_c_11 116.6468396367902
X1045 nt_p_15 nt_c_11 rl_admittance res=22.637692682154487 ind=1.9533517488798835e-06
X1046 nt_n_15 nt_c_11 rl_admittance res=42.23910282158754 ind=1.614574710760359e-05
X1047 nt_n_15 nt_c_11 rl_admittance res=80.38752904923233 ind=6.748332959605176e-05
X1048 nt_p_15 nt_c_11 rl_admittance res=171.8313039832957 ind=0.005840619765153394
X1049 nt_n_15 nt_c_11 rl_admittance res=226.03085108711676 ind=0.8775071639609088
X1050 nt_n_15 nt_c_11 rl_admittance res=1133.947342115307 ind=0.3776963096064935
* Transfer network from port 16 to port 11
R11_16 nt_p_16 nt_c_11 260.5253495067654
X1051 nt_n_16 nt_c_11 rl_admittance res=187.70273079313165 ind=1.6196414652864645e-05
X1052 nt_n_16 nt_c_11 rl_admittance res=223.07021844074174 ind=8.526779911483787e-05
X1053 nt_p_16 nt_c_11 rl_admittance res=145.3572979627057 ind=0.00012202383334361797
X1054 nt_n_16 nt_c_11 rl_admittance res=85.70349740580166 ind=0.0029130986571559688
X1055 nt_n_16 nt_c_11 rl_admittance res=16.297139576480458 ind=0.06326949025609173
X1056 nt_p_16 nt_c_11 rl_admittance res=13.865608639252647 ind=0.004618370729388867

* Port network for port 12
R_ref_12 p12 a12 50.0
H_b_12 a12 0 V_c_12 14.142135623730951
* Differential incident wave a sources for transfer from port 12
H_p_12 nt_p_12 nts_p_12 H_b_12 3.5355339059327378
E_p_12 nts_p_12 0 p12 0 0.07071067811865475
E_n_12 0 nt_n_12 nt_p_12 0 1
* Current sensor on center node for transfer to port 12
V_c_12 nt_c_12 0 0
* Transfer network from port 1 to port 12
R12_1 nt_n_1 nt_c_12 34.746221263150574
X1057 nt_p_1 nt_c_12 rl_admittance res=36.95546541308673 ind=3.1887977281460637e-06
X1058 nt_p_1 nt_c_12 rl_admittance res=83.84323226868591 ind=3.204877789692109e-05
X1059 nt_n_1 nt_c_12 rl_admittance res=112.90233061646438 ind=9.477869613938621e-05
X1060 nt_n_1 nt_c_12 rl_admittance res=41.18713436907605 ind=0.001399968372988892
X1061 nt_n_1 nt_c_12 rl_admittance res=4.464197927787613 ind=0.01733111052819619
X1062 nt_p_1 nt_c_12 rl_admittance res=4.049656806376211 ind=0.0013488637206802317
* Transfer network from port 2 to port 12
R12_2 nt_n_2 nt_c_12 29.061875243318806
X1063 nt_p_2 nt_c_12 rl_admittance res=10.189067843565525 ind=8.791900204288089e-07
X1064 nt_n_2 nt_c_12 rl_admittance res=24.4879261272941 ind=9.360422831682416e-06
X1065 nt_n_2 nt_c_12 rl_admittance res=49.35568609969487 ind=4.143286989783133e-05
X1066 nt_n_2 nt_c_12 rl_admittance res=21.854330313389298 ind=0.0007428380663105547
X1067 nt_n_2 nt_c_12 rl_admittance res=2.3298986553530465 ind=0.009045237636994939
X1068 nt_p_2 nt_c_12 rl_admittance res=2.117194259201725 ind=0.0007051971716154268
* Transfer network from port 3 to port 12
R12_3 nt_n_3 nt_c_12 14.315787610195743
X1069 nt_p_3 nt_c_12 rl_admittance res=7.252729368697202 ind=6.258204754084882e-07
X1070 nt_n_3 nt_c_12 rl_admittance res=25.831320443187 ind=9.873930539973832e-06
X1071 nt_n_3 nt_c_12 rl_admittance res=39.46524431095641 ind=3.313009021329548e-05
X1072 nt_n_3 nt_c_12 rl_admittance res=14.881776902484443 ind=0.0005058379835475355
X1073 nt_n_3 nt_c_12 rl_admittance res=1.7240274821589947 ind=0.006693097243955095
X1074 nt_p_3 nt_c_12 rl_admittance res=1.5545846632658082 ind=0.0005178026072983579
* Transfer network from port 4 to port 12
R12_4 nt_p_4 nt_c_12 3473.29576565795
X1075 nt_p_4 nt_c_12 rl_admittance res=477.4048720531904 ind=4.119411173401106e-05
X1076 nt_n_4 nt_c_12 rl_admittance res=233.22279992966338 ind=8.914858734800294e-05
X1077 nt_p_4 nt_c_12 rl_admittance res=319.03400008613966 ind=0.0002678211015414383
X1078 nt_n_4 nt_c_12 rl_admittance res=39.27690771086235 ind=0.001335038949087352
X1079 nt_n_4 nt_c_12 rl_admittance res=5.074206576064035 ind=0.019699313613598723
X1080 nt_p_4 nt_c_12 rl_admittance res=4.518628550516501 ind=0.0015050692961005908
* Transfer network from port 5 to port 12
R12_5 nt_n_5 nt_c_12 22.324734639677292
X1081 nt_p_5 nt_c_12 rl_admittance res=8.860328797811553 ind=7.645363419258507e-07
X1082 nt_n_5 nt_c_12 rl_admittance res=22.669450160572303 ind=8.665316848869271e-06
X1083 nt_n_5 nt_c_12 rl_admittance res=47.08730481234236 ind=3.952862027261676e-05
X1084 nt_n_5 nt_c_12 rl_admittance res=21.873043698119723 ind=0.0007434741422885387
X1085 nt_n_5 nt_c_12 rl_admittance res=2.4112988018072623 ind=0.009361252956662569
X1086 nt_p_5 nt_c_12 rl_admittance res=2.184776936262752 ind=0.0007277076769724574
* Transfer network from port 6 to port 12
R12_6 nt_n_6 nt_c_12 14.47762593899421
X1087 nt_p_6 nt_c_12 rl_admittance res=6.913257626683745 ind=5.96528279853593e-07
X1088 nt_n_6 nt_c_12 rl_admittance res=20.276433933494857 ind=7.750594891114109e-06
X1089 nt_n_6 nt_c_12 rl_admittance res=44.26946299790151 ind=3.716311221231815e-05
X1090 nt_n_6 nt_c_12 rl_admittance res=17.075764813353754 ind=0.0005804125742052227
X1091 nt_n_6 nt_c_12 rl_admittance res=2.1710467726960325 ind=0.008428535694008924
X1092 nt_p_6 nt_c_12 rl_admittance res=1.9398662033085479 ind=0.0006461325662206056
* Transfer network from port 7 to port 12
R12_7 nt_p_7 nt_c_12 179.21726095370724
X1093 nt_p_7 nt_c_12 rl_admittance res=397.0060555009937 ind=3.425669231034744e-05
X1094 nt_n_7 nt_c_12 rl_admittance res=118.48875364887844 ind=4.5291905455250176e-05
X1095 nt_p_7 nt_c_12 rl_admittance res=3997.4825273536385 ind=0.0033557870746673954
X1096 nt_p_7 nt_c_12 rl_admittance res=494.0368572567377 ind=0.01679252479797555
X1097 nt_p_7 nt_c_12 rl_admittance res=53.161398936280484 ind=0.20638558050108974
X1098 nt_n_7 nt_c_12 rl_admittance res=48.20617015572014 ind=0.016056559146841533
* Transfer network from port 8 to port 12
R12_8 nt_p_8 nt_c_12 215.72815618774936
X1099 nt_n_8 nt_c_12 rl_admittance res=136.04391182491617 ind=1.1738900108717675e-05
X1100 nt_p_8 nt_c_12 rl_admittance res=1418.9169452298936 ind=0.0005423759652552733
X1101 nt_p_8 nt_c_12 rl_admittance res=597.0467212154269 ind=0.0005012058605178319
X1102 nt_p_8 nt_c_12 rl_admittance res=195.50933470338754 ind=0.006645446190943201
X1103 nt_p_8 nt_c_12 rl_admittance res=23.995968532419003 ind=0.09315823124190498
X1104 nt_n_8 nt_c_12 rl_admittance res=21.526974404060137 ind=0.007170226065559383
* Transfer network from port 9 to port 12
R12_9 nt_n_9 nt_c_12 38.40645700682807
X1105 nt_p_9 nt_c_12 rl_admittance res=44.49931481670726 ind=3.839738247250514e-06
X1106 nt_p_9 nt_c_12 rl_admittance res=83.77381437028053 ind=3.202224315168446e-05
X1107 nt_n_9 nt_c_12 rl_admittance res=170.47399584794593 ind=0.0001431086760026835
X1108 nt_n_9 nt_c_12 rl_admittance res=20.861742251597214 ind=0.0007090995721132359
X1109 nt_n_9 nt_c_12 rl_admittance res=2.635350483361616 ind=0.010231076499403895
X1110 nt_p_9 nt_c_12 rl_admittance res=2.3535779050001935 ind=0.0007839320716883539
* Transfer network from port 10 to port 12
R12_10 nt_n_10 nt_c_12 3.725010999427927
X1111 nt_p_10 nt_c_12 rl_admittance res=1.9037181429316432 ind=1.6426723412502733e-07
X1112 nt_n_10 nt_c_12 rl_admittance res=10.857976365932691 ind=4.150422920798605e-06
X1113 nt_n_10 nt_c_12 rl_admittance res=6.409860404139348 ind=5.380918252286398e-06
X1114 nt_n_10 nt_c_12 rl_admittance res=4.2347832740548785 ind=0.00014394210087581233
X1115 nt_n_10 nt_c_12 rl_admittance res=0.29758564986108016 ind=0.0011553004308443471
X1116 nt_p_10 nt_c_12 rl_admittance res=0.27872301153141166 ind=9.283733816196686e-05
* Transfer network from port 11 to port 12
R12_11 nt_n_11 nt_c_12 8.664604329431024
X1117 nt_p_11 nt_c_12 rl_admittance res=6.808326461143266 ind=5.874740233709049e-07
X1118 nt_n_11 nt_c_12 rl_admittance res=100.20223394020591 ind=3.8301948212513964e-05
X1119 nt_n_11 nt_c_12 rl_admittance res=67.70288619581889 ind=5.6834887672170095e-05
X1120 nt_n_11 nt_c_12 rl_admittance res=8.800760932064708 ind=0.00029914164099693907
X1121 nt_n_11 nt_c_12 rl_admittance res=1.9015484744605915 ind=0.00738227724637017
X1122 nt_p_11 nt_c_12 rl_admittance res=1.5802862545519394 ind=0.0005263633189110132
* Transfer network from port 12 to port 12
R12_12 nt_p_12 nt_c_12 1.2585217216533362
X1123 nt_p_12 nt_c_12 rl_admittance res=4.756837051316373 ind=4.104559640325122e-07
X1124 nt_n_12 nt_c_12 rl_admittance res=0.509983952403858 ind=1.9493955539795635e-07
X1125 nt_n_12 nt_c_12 rl_admittance res=37.504448986678184 ind=3.1484051347520344e-05
X1126 nt_p_12 nt_c_12 rl_admittance res=10.547074518349538 ind=0.00035849958923902777
X1127 nt_p_12 nt_c_12 rl_admittance res=0.4638175013822969 ind=0.0018006532217876186
X1128 nt_n_12 nt_c_12 rl_admittance res=0.44456259213184024 ind=0.0001480753507689942
* Transfer network from port 13 to port 12
R12_13 nt_n_13 nt_c_12 12.556224408276842
X1129 nt_p_13 nt_c_12 rl_admittance res=8.011604854110162 ind=6.913020055903174e-07
X1130 nt_n_13 nt_c_12 rl_admittance res=749.6348605766548 ind=0.00028654526430254906
X1131 nt_n_13 nt_c_12 rl_admittance res=23.897631500524305 ind=2.0061466774618713e-05
X1132 nt_n_13 nt_c_12 rl_admittance res=25.81120370116162 ind=0.0008773338908844005
X1133 nt_n_13 nt_c_12 rl_admittance res=2.306168156902193 ind=0.008953110025676246
X1134 nt_p_13 nt_c_12 rl_admittance res=2.126010607742237 ind=0.0007081337297643654
* Transfer network from port 14 to port 12
R12_14 nt_n_14 nt_c_12 21.540314798281393
X1135 nt_p_14 nt_c_12 rl_admittance res=20.174062392851376 ind=1.7407710498761686e-06
X1136 nt_p_14 nt_c_12 rl_admittance res=16.821203436191215 ind=6.42984529935355e-06
X1137 nt_n_14 nt_c_12 rl_admittance res=18.584209571631046 ind=1.5600981329285607e-05
X1138 nt_n_14 nt_c_12 rl_admittance res=5.393368286089146 ind=0.00018332290265076515
X1139 nt_n_14 nt_c_12 rl_admittance res=0.5803272711947403 ind=0.002252972704681796
X1140 nt_p_14 nt_c_12 rl_admittance res=0.5263726221538485 ind=0.0001753247170142276
* Transfer network from port 15 to port 12
R12_15 nt_n_15 nt_c_12 196.67558621106403
X1141 nt_p_15 nt_c_12 rl_admittance res=119.87301015905771 ind=1.0343552115727651e-05
X1142 nt_n_15 nt_c_12 rl_admittance res=1065.8164198361276 ind=0.00040740454290640645
X1143 nt_n_15 nt_c_12 rl_admittance res=499.597269053418 ind=0.00041939947118129666
X1144 nt_n_15 nt_c_12 rl_admittance res=194.6480838242199 ind=0.006616171903947676
X1145 nt_n_15 nt_c_12 rl_admittance res=21.97857661419441 ind=0.08532622135367683
X1146 nt_p_15 nt_c_12 rl_admittance res=19.87321769228546 ind=0.006619391133613531
* Transfer network from port 16 to port 12
R12_16 nt_p_16 nt_c_12 337.31410583952135
X1147 nt_p_16 nt_c_12 rl_admittance res=157.09268920710753 ind=1.3555148199394281e-05
X1148 nt_n_16 nt_c_12 rl_admittance res=112.96226504851599 ind=4.317942480642108e-05
X1149 nt_n_16 nt_c_12 rl_admittance res=1581.0380998362912 ind=0.0013272421289355048
X1150 nt_p_16 nt_c_12 rl_admittance res=358.90798467096835 ind=0.012199436427162376
X1151 nt_p_16 nt_c_12 rl_admittance res=57.24596053941116 ind=0.22224284976830752
X1152 nt_n_16 nt_c_12 rl_admittance res=49.75130653948758 ind=0.016571214711798392

* Port network for port 13
R_ref_13 p13 a13 50.0
H_b_13 a13 0 V_c_13 14.142135623730951
* Differential incident wave a sources for transfer from port 13
H_p_13 nt_p_13 nts_p_13 H_b_13 3.5355339059327378
E_p_13 nts_p_13 0 p13 0 0.07071067811865475
E_n_13 0 nt_n_13 nt_p_13 0 1
* Current sensor on center node for transfer to port 13
V_c_13 nt_c_13 0 0
* Transfer network from port 1 to port 13
R13_1 nt_n_1 nt_c_13 16.340921720129153
X1153 nt_p_1 nt_c_13 rl_admittance res=9.306893100795353 ind=8.030692955474172e-07
X1154 nt_n_1 nt_c_13 rl_admittance res=190.9546692388436 ind=7.299174444043228e-05
X1155 nt_n_1 nt_c_13 rl_admittance res=22.230701903401044 ind=1.866212087175871e-05
X1156 nt_p_1 nt_c_13 rl_admittance res=22.147150097941136 ind=0.0007527911364533949
X1157 nt_p_1 nt_c_13 rl_admittance res=9.309946742725783 ind=0.03614349511822923
X1158 nt_n_1 nt_c_13 rl_admittance res=6.729678229740318 ind=0.0022415279244541973
* Transfer network from port 2 to port 13
R13_2 nt_n_2 nt_c_13 11.4226846959968
X1159 nt_p_2 nt_c_13 rl_admittance res=4.239061442505971 ind=3.657783590664177e-07
X1160 nt_n_2 nt_c_13 rl_admittance res=11.85836712774157 ind=4.532818738180741e-06
X1161 nt_n_2 nt_c_13 rl_admittance res=14.535221252907872 ind=1.2201956424867692e-05
X1162 nt_p_2 nt_c_13 rl_admittance res=16.352164105264247 ind=0.0005558170755983018
X1163 nt_p_2 nt_c_13 rl_admittance res=4.069601788639403 ind=0.015799191600720162
X1164 nt_n_2 nt_c_13 rl_admittance res=3.3100869714862244 ind=0.0011025270638005975
* Transfer network from port 3 to port 13
R13_3 nt_n_3 nt_c_13 7.5112895963681705
X1165 nt_p_3 nt_c_13 rl_admittance res=2.790975394636015 ind=2.408265164095392e-07
X1166 nt_n_3 nt_c_13 rl_admittance res=7.31877135461348 ind=2.7975743691594194e-06
X1167 nt_n_3 nt_c_13 rl_admittance res=10.589862459885152 ind=8.889925927684798e-06
X1168 nt_p_3 nt_c_13 rl_admittance res=13.124229815277195 ind=0.00044609820378814806
X1169 nt_p_3 nt_c_13 rl_admittance res=3.047610199139289 ind=0.011831569760688686
X1170 nt_n_3 nt_c_13 rl_admittance res=2.509911820512994 ind=0.0008360039279046842
* Transfer network from port 4 to port 13
R13_4 nt_p_4 nt_c_13 562.0259763529515
X1171 nt_p_4 nt_c_13 rl_admittance res=223.36122147772502 ind=1.9273299568617393e-05
X1172 nt_n_4 nt_c_13 rl_admittance res=143.8753828250186 ind=5.4995854337019164e-05
X1173 nt_p_4 nt_c_13 rl_admittance res=284.2244211698351 ind=0.00023859932653613744
X1174 nt_n_4 nt_c_13 rl_admittance res=18.263468616424955 ind=0.00062078313618408
X1175 nt_n_4 nt_c_13 rl_admittance res=2.0489018514689863 ind=0.00795433917215066
X1176 nt_p_4 nt_c_13 rl_admittance res=1.8518647079524497 ind=0.0006168209405380159
* Transfer network from port 5 to port 13
R13_5 nt_n_5 nt_c_13 66.11968133022698
X1177 nt_p_5 nt_c_13 rl_admittance res=3.80849687853029 ind=3.286259842260876e-07
X1178 nt_n_5 nt_c_13 rl_admittance res=4.891941610995699 ind=1.8699273147424035e-06
X1179 nt_n_5 nt_c_13 rl_admittance res=23.66104896326002 ind=1.986286162369912e-05
X1180 nt_p_5 nt_c_13 rl_admittance res=592.8232511796205 ind=0.02015031672237547
X1181 nt_p_5 nt_c_13 rl_admittance res=10.958605981466388 ind=0.04254399436851798
X1182 nt_n_5 nt_c_13 rl_admittance res=10.671880259108935 ind=0.003554600501032757
* Transfer network from port 6 to port 13
R13_6 nt_n_6 nt_c_13 7.608688636251869
X1183 nt_p_6 nt_c_13 rl_admittance res=2.587765813591 ind=2.2329205315408826e-07
X1184 nt_n_6 nt_c_13 rl_admittance res=5.482672508744638 ind=2.0957321033523413e-06
X1185 nt_n_6 nt_c_13 rl_admittance res=13.13606446133685 ind=1.102739912675351e-05
X1186 nt_p_6 nt_c_13 rl_admittance res=18.93875329079365 ind=0.000643736352069623
X1187 nt_p_6 nt_c_13 rl_admittance res=3.07821491510179 ind=0.01195038476925463
X1188 nt_n_6 nt_c_13 rl_admittance res=2.6727162910610116 ind=0.0008902310030338681
* Transfer network from port 7 to port 13
R13_7 nt_p_7 nt_c_13 604.7940803433156
X1189 nt_n_7 nt_c_13 rl_admittance res=170.3045307342261 ind=1.4695166049944268e-05
X1190 nt_p_7 nt_c_13 rl_admittance res=489.5058264105562 ind=0.00018711186443297418
X1191 nt_p_7 nt_c_13 rl_admittance res=472.8328738397693 ind=0.0003969314276302194
X1192 nt_p_7 nt_c_13 rl_admittance res=628.533335062691 ind=0.021364117798825563
X1193 nt_p_7 nt_c_13 rl_admittance res=33.057785874207276 ind=0.12833842720931132
X1194 nt_n_7 nt_c_13 rl_admittance res=31.46468626263596 ind=0.010480289024845461
* Transfer network from port 8 to port 13
R13_8 nt_p_8 nt_c_13 101.41839962165247
X1195 nt_n_8 nt_c_13 rl_admittance res=43.27905491365133 ind=3.7344449715978527e-06
X1196 nt_p_8 nt_c_13 rl_admittance res=222.24095654231877 ind=8.495081669798915e-05
X1197 nt_p_8 nt_c_13 rl_admittance res=104.35990325791275 ind=8.760754101364006e-05
X1198 nt_n_8 nt_c_13 rl_admittance res=98.04426832024664 ind=0.0033325667566772555
X1199 nt_n_8 nt_c_13 rl_admittance res=23.858033386970305 ind=0.09262273319944275
X1200 nt_p_8 nt_c_13 rl_admittance res=19.501467246377757 ind=0.006495568124996583
* Transfer network from port 9 to port 13
R13_9 nt_n_9 nt_c_13 26.473335567977948
X1201 nt_p_9 nt_c_13 rl_admittance res=15.266798033197707 ind=1.3173350772382923e-06
X1202 nt_p_9 nt_c_13 rl_admittance res=32.55908882645621 ind=1.2445596121357343e-05
X1203 nt_n_9 nt_c_13 rl_admittance res=15.654671621260828 ind=1.3141707143262307e-05
X1204 nt_p_9 nt_c_13 rl_admittance res=19.564634937758044 ind=0.0006650103378519947
X1205 nt_n_9 nt_c_13 rl_admittance res=35.49608611390727 ind=0.13780450636591143
X1206 nt_n_9 nt_c_13 rl_admittance res=57.13433202159332 ind=0.01903036018950655
* Transfer network from port 10 to port 13
R13_10 nt_n_10 nt_c_13 8.912764118947624
X1207 nt_p_10 nt_c_13 rl_admittance res=5.849145530249447 ind=5.047086207673671e-07
X1208 nt_p_10 nt_c_13 rl_admittance res=303.8364927075862 ind=0.00011614042073854713
X1209 nt_n_10 nt_c_13 rl_admittance res=18.02148740620602 ind=1.5128590078932285e-05
X1210 nt_n_10 nt_c_13 rl_admittance res=7.698393192032006 ind=0.0002616716884234057
X1211 nt_n_10 nt_c_13 rl_admittance res=0.7626363011488628 ind=0.002960741042809444
X1212 nt_p_10 nt_c_13 rl_admittance res=0.6970729737054381 ind=0.00023218176004878013
* Transfer network from port 11 to port 13
R13_11 nt_n_11 nt_c_13 4.942423249070729
X1213 nt_p_11 nt_c_13 rl_admittance res=2.718348478897979 ind=2.345597155096189e-07
X1214 nt_p_11 nt_c_13 rl_admittance res=16.060449665243876 ind=6.139049871033184e-06
X1215 nt_n_11 nt_c_13 rl_admittance res=4.34645527327504 ind=3.6487410080894602e-06
X1216 nt_n_11 nt_c_13 rl_admittance res=21.719240821227878 ind=0.0007382463164972656
X1217 nt_n_11 nt_c_13 rl_admittance res=0.4886763272157343 ind=0.00189716127655794
X1218 nt_p_11 nt_c_13 rl_admittance res=0.47740571274154914 ind=0.0001590147700784551
* Transfer network from port 12 to port 13
R13_12 nt_n_12 nt_c_13 12.560126395464168
X1219 nt_p_12 nt_c_13 rl_admittance res=8.016398902867714 ind=6.917156724624789e-07
X1220 nt_n_12 nt_c_13 rl_admittance res=820.7911667761033 ind=0.0003137445097472306
X1221 nt_n_12 nt_c_13 rl_admittance res=23.85399500983773 ind=2.0024835026905535e-05
X1222 nt_n_12 nt_c_13 rl_admittance res=26.02072631324356 ind=0.0008844556543873493
X1223 nt_n_12 nt_c_13 rl_admittance res=2.315519085595139 ind=0.008989412622769883
X1224 nt_p_12 nt_c_13 rl_admittance res=2.1353273757921505 ind=0.0007112369681416852
* Transfer network from port 13 to port 13
R13_13 nt_p_13 nt_c_13 1.0833634035772979
X1225 nt_n_13 nt_c_13 rl_admittance res=2.645774131167664 ind=2.2829745057594123e-07
X1226 nt_n_13 nt_c_13 rl_admittance res=0.55964484341693 ind=2.139222546949105e-07
X1227 nt_p_13 nt_c_13 rl_admittance res=3.276401000459379 ind=2.7504570823096534e-06
X1228 nt_n_13 nt_c_13 rl_admittance res=1.6188348459196908 ind=5.5024891148569455e-05
X1229 nt_n_13 nt_c_13 rl_admittance res=1.3643865896509408 ind=0.005296883151448411
X1230 nt_p_13 nt_c_13 rl_admittance res=0.7675310265325164 ind=0.0002556499984285309
* Transfer network from port 14 to port 13
R13_14 nt_n_14 nt_c_13 4.768495713152491
X1231 nt_p_14 nt_c_13 rl_admittance res=3.2104311758950086 ind=2.770203412575075e-07
X1232 nt_p_14 nt_c_13 rl_admittance res=10.265116447045038 ind=3.923804321416274e-06
X1233 nt_n_14 nt_c_13 rl_admittance res=5.234566065838255 ind=4.394287911212322e-06
X1234 nt_n_14 nt_c_13 rl_admittance res=5.1163069505019765 ind=0.00017390546895109694
X1235 nt_n_14 nt_c_13 rl_admittance res=0.4443273078393436 ind=0.0017249875134178598
X1236 nt_p_14 nt_c_13 rl_admittance res=0.4101904523816044 ind=0.00013662664424200048
* Transfer network from port 15 to port 13
R13_15 nt_n_15 nt_c_13 184.7323991999749
X1237 nt_p_15 nt_c_13 rl_admittance res=39.93282258171008 ind=3.4457066770406282e-06
X1238 nt_n_15 nt_c_13 rl_admittance res=81.58900154554935 ind=3.118710620536821e-05
X1239 nt_n_15 nt_c_13 rl_admittance res=126.95266373894073 ind=0.00010657360104879951
X1240 nt_p_15 nt_c_13 rl_admittance res=152.6056545792207 ind=0.005187131691069605
X1241 nt_p_15 nt_c_13 rl_admittance res=35.58139179500535 ind=0.13813568392831105
X1242 nt_n_15 nt_c_13 rl_admittance res=29.27992623751663 ind=0.00975258698065349
* Transfer network from port 16 to port 13
R13_16 nt_p_16 nt_c_13 583.6929920898647
X1243 nt_n_16 nt_c_13 rl_admittance res=253.51363063465908 ind=2.187507802663441e-05
X1244 nt_n_16 nt_c_13 rl_admittance res=3054.2961059680056 ind=0.0011674938439623895
X1245 nt_p_16 nt_c_13 rl_admittance res=379.25463932321236 ind=0.0003183748291430346
X1246 nt_n_16 nt_c_13 rl_admittance res=5257.167998905923 ind=0.1786933964379785
X1247 nt_p_16 nt_c_13 rl_admittance res=57.35676743964221 ind=0.2226730293137165
X1248 nt_n_16 nt_c_13 rl_admittance res=57.72052242481044 ind=0.019225609072588575

* Port network for port 14
R_ref_14 p14 a14 50.0
H_b_14 a14 0 V_c_14 14.142135623730951
* Differential incident wave a sources for transfer from port 14
H_p_14 nt_p_14 nts_p_14 H_b_14 3.5355339059327378
E_p_14 nts_p_14 0 p14 0 0.07071067811865475
E_n_14 0 nt_n_14 nt_p_14 0 1
* Current sensor on center node for transfer to port 14
V_c_14 nt_c_14 0 0
* Transfer network from port 1 to port 14
R14_1 nt_n_1 nt_c_14 14.540363199534857
X1249 nt_p_1 nt_c_14 rl_admittance res=8.981058107521708 ind=7.749537820587534e-07
X1250 nt_p_1 nt_c_14 rl_admittance res=91.59267682955662 ind=3.501097557031168e-05
X1251 nt_n_1 nt_c_14 rl_admittance res=19.686294982142233 ind=1.652615459782802e-05
X1252 nt_n_1 nt_c_14 rl_admittance res=18.4146430582096 ind=0.0006259216203380457
X1253 nt_n_1 nt_c_14 rl_admittance res=1.4301475701286601 ind=0.005552183395644063
X1254 nt_p_1 nt_c_14 rl_admittance res=1.331840066405304 ind=0.0004436106152239643
* Transfer network from port 2 to port 14
R14_2 nt_n_2 nt_c_14 7.242167421676161
X1255 nt_p_2 nt_c_14 rl_admittance res=4.147592800906233 ind=3.5788575121343793e-07
X1256 nt_p_2 nt_c_14 rl_admittance res=451.14785996353055 ind=0.00017244966792677615
X1257 nt_n_2 nt_c_14 rl_admittance res=10.090893531805753 ind=8.471053933110257e-06
X1258 nt_n_2 nt_c_14 rl_admittance res=8.473242706225134 ind=0.0002880091559436187
X1259 nt_n_2 nt_c_14 rl_admittance res=0.6864331984553291 ind=0.002664901920813429
X1260 nt_p_2 nt_c_14 rl_admittance res=0.6374769013992216 ind=0.00021233144095449998
* Transfer network from port 3 to port 14
R14_3 nt_n_3 nt_c_14 5.075373106598556
X1261 nt_p_3 nt_c_14 rl_admittance res=2.2684804090115676 ind=1.9574168783268316e-07
X1262 nt_n_3 nt_c_14 rl_admittance res=11.1023605381343 ind=4.243837903075444e-06
X1263 nt_n_3 nt_c_14 rl_admittance res=6.900844441195517 ind=5.793087129610261e-06
X1264 nt_n_3 nt_c_14 rl_admittance res=6.115171592180823 ind=0.0002078573067924106
X1265 nt_n_3 nt_c_14 rl_admittance res=0.527256288683986 ind=0.002046938142905617
X1266 nt_p_3 nt_c_14 rl_admittance res=0.48748958530274256 ind=0.00016237351639007848
* Transfer network from port 4 to port 14
R14_4 nt_p_4 nt_c_14 1348.3715623673531
X1267 nt_p_4 nt_c_14 rl_admittance res=181.835820818317 ind=1.5690173181141727e-05
X1268 nt_n_4 nt_c_14 rl_admittance res=87.38253858818037 ind=3.340166517325062e-05
X1269 nt_p_4 nt_c_14 rl_admittance res=81.48202524270933 ind=6.840213190580803e-05
X1270 nt_n_4 nt_c_14 rl_admittance res=7.165427683856979 ind=0.00024355596207417953
X1271 nt_n_4 nt_c_14 rl_admittance res=0.8151964449895993 ind=0.0031647924036623293
X1272 nt_p_4 nt_c_14 rl_admittance res=0.7357337160771505 ind=0.00024505891860642886
* Transfer network from port 5 to port 14
R14_5 nt_n_5 nt_c_14 7.823577605451835
X1273 nt_p_5 nt_c_14 rl_admittance res=3.194706689318662 ind=2.7566351334286947e-07
X1274 nt_n_5 nt_c_14 rl_admittance res=17.15197417644752 ind=6.556281240602845e-06
X1275 nt_n_5 nt_c_14 rl_admittance res=8.288287877117714 ind=6.9578113572311165e-06
X1276 nt_n_5 nt_c_14 rl_admittance res=8.437437185156918 ind=0.00028679211091628783
X1277 nt_n_5 nt_c_14 rl_admittance res=0.6907301480009341 ind=0.0026815837321295033
X1278 nt_p_5 nt_c_14 rl_admittance res=0.6410178956283418 ind=0.00021351087883755168
* Transfer network from port 6 to port 14
R14_6 nt_n_6 nt_c_14 5.414728302179013
X1279 nt_p_6 nt_c_14 rl_admittance res=1.9107213202657702 ind=1.648715213589519e-07
X1280 nt_n_6 nt_c_14 rl_admittance res=5.1043983099364 ind=1.9511381337056246e-06
X1281 nt_n_6 nt_c_14 rl_admittance res=7.468665064060158 ind=6.269758408071157e-06
X1282 nt_n_6 nt_c_14 rl_admittance res=6.208147607920204 ind=0.00021101760146878364
X1283 nt_n_6 nt_c_14 rl_admittance res=0.5718960318937041 ind=0.00222024056722293
X1284 nt_p_6 nt_c_14 rl_admittance res=0.5261025474051244 ind=0.00017523476024805122
* Transfer network from port 7 to port 14
R14_7 nt_p_7 nt_c_14 544.0915521659688
X1285 nt_n_7 nt_c_14 rl_admittance res=58.61107507858343 ind=5.057407908833975e-06
X1286 nt_p_7 nt_c_14 rl_admittance res=109.67344913202457 ind=4.192228659741552e-05
X1287 nt_p_7 nt_c_14 rl_admittance res=164.5126172966239 ind=0.000138104247102035
X1288 nt_p_7 nt_c_14 rl_admittance res=1472.8806989930968 ind=0.050063847057159674
X1289 nt_p_7 nt_c_14 rl_admittance res=32.99938182729383 ind=0.12811168838439266
X1290 nt_n_7 nt_c_14 rl_admittance res=32.30462610865816 ind=0.010760057024955798
* Transfer network from port 8 to port 14
R14_8 nt_p_8 nt_c_14 70.01605554952133
X1291 nt_n_8 nt_c_14 rl_admittance res=47.162304566683325 ind=4.069521191934869e-06
X1292 nt_n_8 nt_c_14 rl_admittance res=188.57067252715075 ind=7.208047016041422e-05
X1293 nt_p_8 nt_c_14 rl_admittance res=86.76267801205486 ind=7.283510845740475e-05
X1294 nt_p_8 nt_c_14 rl_admittance res=74.86663832046342 ind=0.0025447491661216596
X1295 nt_p_8 nt_c_14 rl_admittance res=6.600438643451615 ind=0.025624520577860806
X1296 nt_n_8 nt_c_14 rl_admittance res=6.091474033020952 ind=0.002028954235250409
* Transfer network from port 9 to port 14
R14_9 nt_n_9 nt_c_14 16.0247084301923
X1297 nt_p_9 nt_c_14 rl_admittance res=11.067933513793154 ind=9.55025213443994e-07
X1298 nt_p_9 nt_c_14 rl_admittance res=29.336484774183834 ind=1.1213767162401892e-05
X1299 nt_n_9 nt_c_14 rl_admittance res=16.475732134832125 ind=1.3830967006215694e-05
X1300 nt_n_9 nt_c_14 rl_admittance res=21.00319453358627 ind=0.000713907595883408
X1301 nt_n_9 nt_c_14 rl_admittance res=1.4917116335574176 ind=0.005791190179193522
X1302 nt_p_9 nt_c_14 rl_admittance res=1.3953935810700557 ind=0.0004647790831588342
* Transfer network from port 10 to port 14
R14_10 nt_n_10 nt_c_14 11.126548996156195
X1303 nt_p_10 nt_c_14 rl_admittance res=12.632941424017954 ind=1.0900659608103693e-06
X1304 nt_p_10 nt_c_14 rl_admittance res=13.501092368404468 ind=5.16074462986102e-06
X1305 nt_n_10 nt_c_14 rl_admittance res=18.321624870736848 ind=1.538054800925569e-05
X1306 nt_n_10 nt_c_14 rl_admittance res=6.265647302753542 ind=0.00021297204077261694
X1307 nt_n_10 nt_c_14 rl_admittance res=0.983596079425552 ind=0.0038185610592030394
X1308 nt_p_10 nt_c_14 rl_admittance res=0.8565259649537168 ind=0.00028529252111626123
* Transfer network from port 11 to port 14
R14_11 nt_n_11 nt_c_14 3.2811495353743
X1309 nt_p_11 nt_c_14 rl_admittance res=2.680355524305895 ind=2.3128139534954077e-07
X1310 nt_p_11 nt_c_14 rl_admittance res=5.992785617536668 ind=2.29072102832118e-06
X1311 nt_n_11 nt_c_14 rl_admittance res=4.50581154025299 ind=3.7825166274530488e-06
X1312 nt_n_11 nt_c_14 rl_admittance res=3.963279806270113 ind=0.0001347135814879507
X1313 nt_n_11 nt_c_14 rl_admittance res=0.6800868952385232 ind=0.002640264016250264
X1314 nt_p_11 nt_c_14 rl_admittance res=0.5849760630502726 ind=0.00019484440945032565
* Transfer network from port 12 to port 14
R14_12 nt_n_12 nt_c_14 21.513960365804525
X1315 nt_p_12 nt_c_14 rl_admittance res=20.12731458474947 ind=1.736737294581657e-06
X1316 nt_p_12 nt_c_14 rl_admittance res=16.81696277553374 ind=6.428224321871289e-06
X1317 nt_n_12 nt_c_14 rl_admittance res=18.55690212388313 ind=1.5578057406649908e-05
X1318 nt_n_12 nt_c_14 rl_admittance res=5.397974824952458 ind=0.00018347948088366168
X1319 nt_n_12 nt_c_14 rl_admittance res=0.5803469317460141 ind=0.0022530490317606323
X1320 nt_p_12 nt_c_14 rl_admittance res=0.5264309985619201 ind=0.0001753441610863444
* Transfer network from port 13 to port 14
R14_13 nt_n_13 nt_c_14 4.76679999518172
X1321 nt_p_13 nt_c_14 rl_admittance res=3.209125841788304 ind=2.7690770713458676e-07
X1322 nt_p_13 nt_c_14 rl_admittance res=10.283386145469322 ind=3.9307878487827665e-06
X1323 nt_n_13 nt_c_14 rl_admittance res=5.238071986464991 ind=4.39723104430759e-06
X1324 nt_n_13 nt_c_14 rl_admittance res=5.11178127685578 ind=0.00017375163936163415
X1325 nt_n_13 nt_c_14 rl_admittance res=0.4441921946971727 ind=0.0017244629710837934
X1326 nt_p_13 nt_c_14 rl_admittance res=0.41004735812060433 ind=0.0001365789822630899
* Transfer network from port 14 to port 14
R14_14 nt_p_14 nt_c_14 1.5896902532847592
X1327 nt_p_14 nt_c_14 rl_admittance res=1.9793009494760279 ind=1.7078909169336113e-07
X1328 nt_n_14 nt_c_14 rl_admittance res=0.6486665082661809 ind=2.4795047006266837e-07
X1329 nt_n_14 nt_c_14 rl_admittance res=1.7714074395767303 ind=1.487052450892521e-06
X1330 nt_n_14 nt_c_14 rl_admittance res=7.843215489026569 ind=0.0002665942604498834
X1331 nt_n_14 nt_c_14 rl_admittance res=2.022463640202728 ind=0.007851699556023602
X1332 nt_p_14 nt_c_14 rl_admittance res=1.6243217268922594 ind=0.0005410306978773871
* Transfer network from port 15 to port 14
R14_15 nt_n_15 nt_c_14 68.30583783635747
X1333 nt_p_15 nt_c_14 rl_admittance res=45.02798177841364 ind=3.885355640715627e-06
X1334 nt_p_15 nt_c_14 rl_admittance res=170.26180878991778 ind=6.508197199208056e-05
X1335 nt_n_15 nt_c_14 rl_admittance res=78.1044148460338 ind=6.556671205472252e-05
X1336 nt_n_15 nt_c_14 rl_admittance res=81.04486042936301 ind=0.0027547495870359684
X1337 nt_n_15 nt_c_14 rl_admittance res=6.5539948545943805 ind=0.025444214406169213
X1338 nt_p_15 nt_c_14 rl_admittance res=6.08719773579351 ind=0.00202752988191265
* Transfer network from port 16 to port 14
R14_16 nt_p_16 nt_c_14 249.056060411088
X1339 nt_n_16 nt_c_14 rl_admittance res=54.15372513487299 ind=4.672793962962182e-06
X1340 nt_p_16 nt_c_14 rl_admittance res=110.34708778107753 ind=4.217978257964454e-05
X1341 nt_p_16 nt_c_14 rl_admittance res=186.32091869417513 ind=0.00015641177326370696
X1342 nt_p_16 nt_c_14 rl_admittance res=918.7622227783752 ind=0.03122912224630097
X1343 nt_p_16 nt_c_14 rl_admittance res=30.122599381965912 ind=0.11694331383379082
X1344 nt_n_16 nt_c_14 rl_admittance res=29.18496568820293 ind=0.009720957426350655

* Port network for port 15
R_ref_15 p15 a15 50.0
H_b_15 a15 0 V_c_15 14.142135623730951
* Differential incident wave a sources for transfer from port 15
H_p_15 nt_p_15 nts_p_15 H_b_15 3.5355339059327378
E_p_15 nts_p_15 0 p15 0 0.07071067811865475
E_n_15 0 nt_n_15 nt_p_15 0 1
* Current sensor on center node for transfer to port 15
V_c_15 nt_c_15 0 0
* Transfer network from port 1 to port 15
R15_1 nt_p_1 nt_c_15 38.69537240924798
X1345 nt_n_1 nt_c_15 rl_admittance res=69.65522232089367 ind=6.010380662442382e-06
X1346 nt_n_1 nt_c_15 rl_admittance res=73.00501197755749 ind=2.790590666558369e-05
X1347 nt_p_1 nt_c_15 rl_admittance res=293.9204632774792 ind=0.0002467389125274746
X1348 nt_n_1 nt_c_15 rl_admittance res=63.65056847190319 ind=0.0021635101385041413
X1349 nt_n_1 nt_c_15 rl_admittance res=9.194259372210654 ind=0.03569436839097685
X1350 nt_p_1 nt_c_15 rl_admittance res=8.11140210009978 ind=0.002701753886760745
* Transfer network from port 2 to port 15
R15_2 nt_p_2 nt_c_15 18.59450417603047
X1351 nt_n_2 nt_c_15 rl_admittance res=29.494684892676243 ind=2.5450250220592268e-06
X1352 nt_n_2 nt_c_15 rl_admittance res=42.819057333443645 ind=1.6367432660961435e-05
X1353 nt_p_2 nt_c_15 rl_admittance res=176.07470971303388 ind=0.00014781033587705822
X1354 nt_n_2 nt_c_15 rl_admittance res=33.99321803037448 ind=0.001155444069310414
X1355 nt_n_2 nt_c_15 rl_admittance res=4.696146176122018 ind=0.01823159047862197
X1356 nt_p_2 nt_c_15 rl_admittance res=4.163926180741572 ind=0.0013869246776540619
* Transfer network from port 3 to port 15
R15_3 nt_p_3 nt_c_15 15.402631497275504
X1357 nt_n_3 nt_c_15 rl_admittance res=25.638248616789603 ind=2.2122624631838996e-06
X1358 nt_n_3 nt_c_15 rl_admittance res=33.16381383768811 ind=1.2676750110167987e-05
X1359 nt_p_3 nt_c_15 rl_admittance res=139.56788613023193 ind=0.00011716376622277342
X1360 nt_n_3 nt_c_15 rl_admittance res=25.292026865628824 ind=0.0008596868474358015
X1361 nt_n_3 nt_c_15 rl_admittance res=3.496880561598475 ind=0.013575747423680817
X1362 nt_p_3 nt_c_15 rl_admittance res=3.100045201256436 ind=0.0010325661418665885
* Transfer network from port 4 to port 15
R15_4 nt_p_4 nt_c_15 1269.8476950003355
X1363 nt_n_4 nt_c_15 rl_admittance res=8500.427237423486 ind=0.0007334813067559979
X1364 nt_n_4 nt_c_15 rl_admittance res=676.5826342002986 ind=0.00025862131010063246
X1365 nt_p_4 nt_c_15 rl_admittance res=1055.5028860291388 ind=0.0008860683987918702
X1366 nt_n_4 nt_c_15 rl_admittance res=314.74877799572283 ind=0.010698446040998481
X1367 nt_n_4 nt_c_15 rl_admittance res=49.52424970899331 ind=0.19226527573743044
X1368 nt_p_4 nt_c_15 rl_admittance res=43.04750550262995 ind=0.014338305988511452
* Transfer network from port 5 to port 15
R15_5 nt_n_5 nt_c_15 156.3452413000715
X1369 nt_p_5 nt_c_15 rl_admittance res=38.30862522420933 ind=3.3055586154273883e-06
X1370 nt_n_5 nt_c_15 rl_admittance res=45.034250649859516 ind=1.7214182442375472e-05
X1371 nt_p_5 nt_c_15 rl_admittance res=222.99265136095087 ind=0.00018719677998900024
X1372 nt_n_5 nt_c_15 rl_admittance res=36.21027903334668 ind=0.001230802924270678
X1373 nt_n_5 nt_c_15 rl_admittance res=4.8846918906707035 ind=0.018963571154953774
X1374 nt_p_5 nt_c_15 rl_admittance res=4.341203698163113 ind=0.0014459724496444374
* Transfer network from port 6 to port 15
R15_6 nt_n_6 nt_c_15 32.48338337365508
X1375 nt_p_6 nt_c_15 rl_admittance res=17.26963769691129 ind=1.4901552676512927e-06
X1376 nt_n_6 nt_c_15 rl_admittance res=31.538852458938276 ind=1.2055614391643473e-05
X1377 nt_p_6 nt_c_15 rl_admittance res=135.13359108625207 ind=0.00011344128591372243
X1378 nt_n_6 nt_c_15 rl_admittance res=25.847146266246185 ind=0.0008785555940966605
X1379 nt_n_6 nt_c_15 rl_admittance res=3.5971725624475233 ind=0.013965105552492597
X1380 nt_p_6 nt_c_15 rl_admittance res=3.1860139360749806 ind=0.0010612006936456268
* Transfer network from port 7 to port 15
R15_7 nt_n_7 nt_c_15 89.62621112727908
X1381 nt_p_7 nt_c_15 rl_admittance res=87.84320495748202 ind=7.579777693783102e-06
X1382 nt_n_7 nt_c_15 rl_admittance res=4536.840550793469 ind=0.0017341911950647642
X1383 nt_n_7 nt_c_15 rl_admittance res=9792.990316535343 ind=0.008220971599425085
X1384 nt_p_7 nt_c_15 rl_admittance res=704.9521972967026 ind=0.02396162772191788
X1385 nt_p_7 nt_c_15 rl_admittance res=92.76389906129018 ind=0.36013219253797885
X1386 nt_n_7 nt_c_15 rl_admittance res=82.62736127519314 ind=0.027521603752733607
* Transfer network from port 8 to port 15
R15_8 nt_n_8 nt_c_15 12.706269461367498
X1387 nt_p_8 nt_c_15 rl_admittance res=12.433564607827535 ind=1.0728622175641034e-06
X1388 nt_n_8 nt_c_15 rl_admittance res=564.1982048645827 ind=0.00021566276094415167
X1389 nt_n_8 nt_c_15 rl_admittance res=4582.587420034715 ind=0.003846968067391747
X1390 nt_p_8 nt_c_15 rl_admittance res=278.65406783612576 ind=0.009471571352343847
X1391 nt_p_8 nt_c_15 rl_admittance res=38.39578448454794 ind=0.14906184615525844
X1392 nt_n_8 nt_c_15 rl_admittance res=34.04983865299804 ind=0.011341354156660793
* Transfer network from port 9 to port 15
R15_9 nt_n_9 nt_c_15 357.3804467605407
X1393 nt_p_9 nt_c_15 rl_admittance res=51.27396516699876 ind=4.424306440466756e-06
X1394 nt_n_9 nt_c_15 rl_admittance res=50.11492972824877 ind=1.9156253984023863e-05
X1395 nt_p_9 nt_c_15 rl_admittance res=219.11775583487113 ind=0.00018394390165041419
X1396 nt_n_9 nt_c_15 rl_admittance res=61.693690600237616 ind=0.002096995019836635
X1397 nt_n_9 nt_c_15 rl_admittance res=10.610090377822074 ind=0.041190971374182685
X1398 nt_p_9 nt_c_15 rl_admittance res=9.162171450878247 ind=0.0030517451882053955
* Transfer network from port 10 to port 15
R15_10 nt_n_10 nt_c_15 131.81303523384463
X1399 nt_p_10 nt_c_15 rl_admittance res=55.305397412498735 ind=4.772168978305956e-06
X1400 nt_n_10 nt_c_15 rl_admittance res=163.96070622649756 ind=6.267339790569962e-05
X1401 nt_n_10 nt_c_15 rl_admittance res=237.85792089355556 ind=0.00019967580372897038
X1402 nt_n_10 nt_c_15 rl_admittance res=222.44402429055532 ind=0.007560967849245792
X1403 nt_n_10 nt_c_15 rl_admittance res=18.29824880649226 ind=0.07103828675779963
X1404 nt_p_10 nt_c_15 rl_admittance res=16.962411749331686 ind=0.005649856992298443
* Transfer network from port 11 to port 15
R15_11 nt_n_11 nt_c_15 116.18487197670112
X1405 nt_p_11 nt_c_15 rl_admittance res=22.610218435594714 ind=1.9509810625948367e-06
X1406 nt_n_11 nt_c_15 rl_admittance res=42.14232226413012 ind=1.6108753083079907e-05
X1407 nt_n_11 nt_c_15 rl_admittance res=80.70685501381683 ind=6.775139579452188e-05
X1408 nt_p_11 nt_c_15 rl_admittance res=183.13126632110618 ind=0.006224710334483654
X1409 nt_n_11 nt_c_15 rl_admittance res=135.63470523234648 ind=0.526567169705685
X1410 nt_p_11 nt_c_15 rl_admittance res=414.75553022309055 ind=0.13814718491417954
* Transfer network from port 12 to port 15
R15_12 nt_n_12 nt_c_15 195.57658919721663
X1411 nt_p_12 nt_c_15 rl_admittance res=120.11769771625403 ind=1.0364665613224476e-05
X1412 nt_n_12 nt_c_15 rl_admittance res=1143.9521772646567 ind=0.00043727165880682586
X1413 nt_n_12 nt_c_15 rl_admittance res=494.2613115056605 ind=0.0004149200676448933
X1414 nt_n_12 nt_c_15 rl_admittance res=193.92360159443987 ind=0.0065915464420401824
X1415 nt_n_12 nt_c_15 rl_admittance res=22.100907522504844 ind=0.08580113992297814
X1416 nt_p_12 nt_c_15 rl_admittance res=19.964472962944434 ind=0.0066497865300132785
* Transfer network from port 13 to port 15
R15_13 nt_n_13 nt_c_15 184.89879945622243
X1417 nt_p_13 nt_c_15 rl_admittance res=39.884453622848554 ind=3.441533036568066e-06
X1418 nt_n_13 nt_c_15 rl_admittance res=80.99015565996221 ind=3.0958199491464774e-05
X1419 nt_n_13 nt_c_15 rl_admittance res=128.21854977521147 ind=0.00010763628086527179
X1420 nt_p_13 nt_c_15 rl_admittance res=162.91156495104914 ind=0.005537434007470882
X1421 nt_p_13 nt_c_15 rl_admittance res=40.62713023837495 ind=0.15772447727326586
X1422 nt_n_13 nt_c_15 rl_admittance res=33.03600582748272 ind=0.011003665709822735
* Transfer network from port 14 to port 15
R15_14 nt_n_14 nt_c_15 68.21830783034511
X1423 nt_p_14 nt_c_15 rl_admittance res=44.95471862635035 ind=3.8790339405220335e-06
X1424 nt_p_14 nt_c_15 rl_admittance res=172.38381295506355 ind=6.589310055123676e-05
X1425 nt_n_14 nt_c_15 rl_admittance res=78.59869111543767 ind=6.598164467915063e-05
X1426 nt_n_14 nt_c_15 rl_admittance res=77.72459627683179 ind=0.0026418923835738488
X1427 nt_n_14 nt_c_15 rl_admittance res=6.367679409439323 ind=0.02472089218226131
X1428 nt_p_14 nt_c_15 rl_admittance res=5.908590206830401 ind=0.0019680391083539235
* Transfer network from port 15 to port 15
R15_15 nt_n_15 nt_c_15 2.798691986927389
X1429 nt_n_15 nt_c_15 rl_admittance res=1.4514232136147982 ind=1.2523979861756384e-07
X1430 nt_p_15 nt_c_15 rl_admittance res=17.927469703433662 ind=6.852711652836809e-06
X1431 nt_n_15 nt_c_15 rl_admittance res=121.99174959587697 ind=0.00010240903711489559
X1432 nt_n_15 nt_c_15 rl_admittance res=255.34122361785415 ind=0.008679157772473581
X1433 nt_n_15 nt_c_15 rl_admittance res=98.8890838348628 ind=0.38391166110850006
X1434 nt_p_15 nt_c_15 rl_admittance res=72.81029921136074 ind=0.024251726947192874
* Transfer network from port 16 to port 15
R15_16 nt_n_16 nt_c_15 5667.3260177966595
X1435 nt_n_16 nt_c_15 rl_admittance res=2851.540940353675 ind=0.000246052570862638
X1436 nt_p_16 nt_c_15 rl_admittance res=1472.071120662783 ind=0.0005626939601207801
X1437 nt_n_16 nt_c_15 rl_admittance res=3977.3728301353503 ind=0.0033389054844318324
X1438 nt_p_16 nt_c_15 rl_admittance res=713.2294881661837 ind=0.02424297639083629
X1439 nt_p_16 nt_c_15 rl_admittance res=101.27134227969624 ind=0.39316017228161426
X1440 nt_n_16 nt_c_15 rl_admittance res=89.46713241357834 ind=0.0297998015328016

* Port network for port 16
R_ref_16 p16 a16 50.0
H_b_16 a16 0 V_c_16 14.142135623730951
* Differential incident wave a sources for transfer from port 16
H_p_16 nt_p_16 nts_p_16 H_b_16 3.5355339059327378
E_p_16 nts_p_16 0 p16 0 0.07071067811865475
E_n_16 0 nt_n_16 nt_p_16 0 1
* Current sensor on center node for transfer to port 16
V_c_16 nt_c_16 0 0
* Transfer network from port 1 to port 16
R16_1 nt_n_1 nt_c_16 23.879244335160266
X1441 nt_p_1 nt_c_16 rl_admittance res=26.83949450736334 ind=2.3159150656877192e-06
X1442 nt_p_1 nt_c_16 rl_admittance res=136.38463368767907 ind=5.2132542070922175e-05
X1443 nt_n_1 nt_c_16 rl_admittance res=267.6843310252381 ind=0.00022471433258275126
X1444 nt_p_1 nt_c_16 rl_admittance res=82.04312638583727 ind=0.002788681075310248
X1445 nt_p_1 nt_c_16 rl_admittance res=13.091298362582265 ind=0.05082362891377188
X1446 nt_n_1 nt_c_16 rl_admittance res=11.42166057252237 ind=0.0038043380742639648
* Transfer network from port 2 to port 16
R16_2 nt_p_2 nt_c_16 22.740436863766174
X1447 nt_n_2 nt_c_16 rl_admittance res=20.143938241436103 ind=1.7381717097103338e-06
X1448 nt_p_2 nt_c_16 rl_admittance res=130.34971828220588 ind=4.9825717080720146e-05
X1449 nt_n_2 nt_c_16 rl_admittance res=329.2472234871628 ind=0.0002763948483546691
X1450 nt_p_2 nt_c_16 rl_admittance res=74.31565751990338 ind=0.0025260210922528623
X1451 nt_p_2 nt_c_16 rl_admittance res=10.802116155880919 ind=0.04193646251002262
X1452 nt_n_2 nt_c_16 rl_admittance res=9.524098899336622 ind=0.003172296343052691
* Transfer network from port 3 to port 16
R16_3 nt_p_3 nt_c_16 59.95312655073761
X1453 nt_n_3 nt_c_16 rl_admittance res=38.23487174205105 ind=3.299194605835836e-06
X1454 nt_p_3 nt_c_16 rl_admittance res=85.18828919504126 ind=3.256292113215962e-05
X1455 nt_n_3 nt_c_16 rl_admittance res=298.2639531295098 ind=0.00025038516413824585
X1456 nt_p_3 nt_c_16 rl_admittance res=62.85635894369169 ind=0.0021365146157989404
X1457 nt_p_3 nt_c_16 rl_admittance res=8.803694086622315 ind=0.034178098224980295
X1458 nt_n_3 nt_c_16 rl_admittance res=7.787585808417493 ind=0.0025938968339537702
* Transfer network from port 4 to port 16
R16_4 nt_p_4 nt_c_16 168.92122466436743
X1459 nt_n_4 nt_c_16 rl_admittance res=159.96021103910593 ind=1.3802579722744753e-05
X1460 nt_p_4 nt_c_16 rl_admittance res=1873.9144429406408 ind=0.0007162971435449704
X1461 nt_n_4 nt_c_16 rl_admittance res=4103.357252822737 ind=0.003444666271219723
X1462 nt_p_4 nt_c_16 rl_admittance res=1001.0060071326583 ind=0.034024623772072646
X1463 nt_p_4 nt_c_16 rl_admittance res=136.6930626037224 ind=0.530675972424192
X1464 nt_n_4 nt_c_16 rl_admittance res=120.87564475183719 ind=0.04026138009099191
* Transfer network from port 5 to port 16
R16_5 nt_n_5 nt_c_16 202.71581400217508
X1465 nt_p_5 nt_c_16 rl_admittance res=973.1519527249011 ind=8.397092828632503e-05
X1466 nt_p_5 nt_c_16 rl_admittance res=248.75750323738953 ind=9.508667254023885e-05
X1467 nt_n_5 nt_c_16 rl_admittance res=1494.1984744297263 ind=0.0012543424250558164
X1468 nt_p_5 nt_c_16 rl_admittance res=173.04254304473716 ind=0.005881790300664598
X1469 nt_p_5 nt_c_16 rl_admittance res=23.43687203075641 ind=0.09098768158819723
X1470 nt_n_5 nt_c_16 rl_admittance res=20.880299143176348 ind=0.006954830825870389
* Transfer network from port 6 to port 16
R16_6 nt_n_6 nt_c_16 22.947390300148292
X1471 nt_p_6 nt_c_16 rl_admittance res=28.391427296410072 ind=2.449827592471785e-06
X1472 nt_p_6 nt_c_16 rl_admittance res=103.88968530558148 ind=3.971146340672669e-05
X1473 nt_n_6 nt_c_16 rl_admittance res=500.9255606573881 ind=0.0004205145389184264
X1474 nt_p_6 nt_c_16 rl_admittance res=100.35359141075283 ind=0.003411061639587803
X1475 nt_p_6 nt_c_16 rl_admittance res=13.906029755477256 ind=0.05398661587121892
X1476 nt_n_6 nt_c_16 rl_admittance res=12.322970367856156 ind=0.004104547238187503
* Transfer network from port 7 to port 16
R16_7 nt_p_7 nt_c_16 6.097855579465656
X1477 nt_n_7 nt_c_16 rl_admittance res=5.929043885493943 ind=5.116028565952302e-07
X1478 nt_p_7 nt_c_16 rl_admittance res=217.94188783816082 ind=8.33075129472269e-05
X1479 nt_p_7 nt_c_16 rl_admittance res=3875.3038088479634 ind=0.0032532210818068345
X1480 nt_n_7 nt_c_16 rl_admittance res=704.6284653496054 ind=0.023950623934103927
X1481 nt_n_7 nt_c_16 rl_admittance res=119.6314856993349 ind=0.4644387490979848
X1482 nt_p_7 nt_c_16 rl_admittance res=104.15637562163212 ind=0.03469250928433139
* Transfer network from port 8 to port 16
R16_8 nt_p_8 nt_c_16 88.20213713345609
X1483 nt_n_8 nt_c_16 rl_admittance res=88.6113509932816 ind=7.646059157335574e-06
X1484 nt_n_8 nt_c_16 rl_admittance res=5767.972456614255 ind=0.002204786995630051
X1485 nt_p_8 nt_c_16 rl_admittance res=4288.707232268728 ind=0.0036002629651536145
X1486 nt_n_8 nt_c_16 rl_admittance res=497.65189943837373 ind=0.016915401633153263
X1487 nt_n_8 nt_c_16 rl_admittance res=66.71681126907204 ind=0.2590110136013
X1488 nt_p_8 nt_c_16 rl_admittance res=59.220639031238505 ind=0.01972526940529006
* Transfer network from port 9 to port 16
R16_9 nt_n_9 nt_c_16 31.249990277285995
X1489 nt_p_9 nt_c_16 rl_admittance res=252.7885108828272 ind=2.1812509197059972e-05
X1490 nt_p_9 nt_c_16 rl_admittance res=23.042528912505706 ind=8.807924877391567e-06
X1491 nt_n_9 nt_c_16 rl_admittance res=49.92413004191518 ind=4.1910064437375375e-05
X1492 nt_p_9 nt_c_16 rl_admittance res=16.554655480301466 ind=0.0005626998443365896
X1493 nt_p_9 nt_c_16 rl_admittance res=2.6234569852668206 ind=0.010184903024709879
X1494 nt_n_9 nt_c_16 rl_admittance res=2.2888225328522522 ind=0.0007623632878664809
* Transfer network from port 10 to port 16
R16_10 nt_p_10 nt_c_16 116.61215500847871
X1495 nt_p_10 nt_c_16 rl_admittance res=92.665591635792 ind=7.995889776587266e-06
X1496 nt_n_10 nt_c_16 rl_admittance res=47.17049175311182 ind=1.8030753020582736e-05
X1497 nt_p_10 nt_c_16 rl_admittance res=483.16510401685247 ind=0.0004056050776695849
X1498 nt_n_10 nt_c_16 rl_admittance res=399.9610187758162 ind=0.013594846674619967
X1499 nt_n_10 nt_c_16 rl_admittance res=523.7487844251685 ind=2.033321151685469
X1500 nt_p_10 nt_c_16 rl_admittance res=239.65006476327767 ind=0.07982288215359032
* Transfer network from port 11 to port 16
R16_11 nt_p_11 nt_c_16 258.79199803603643
X1501 nt_n_11 nt_c_16 rl_admittance res=187.18356461643697 ind=1.615161705915911e-05
X1502 nt_n_11 nt_c_16 rl_admittance res=226.60051128667433 ind=8.66172410228956e-05
X1503 nt_p_11 nt_c_16 rl_admittance res=147.7157365145378 ind=0.00012400368380061918
X1504 nt_n_11 nt_c_16 rl_admittance res=89.57462765920597 ind=0.0030446800357953026
X1505 nt_n_11 nt_c_16 rl_admittance res=17.53197061565191 ind=0.06806340700658263
X1506 nt_p_11 nt_c_16 rl_admittance res=14.853557203385442 ind=0.004947437620676705
* Transfer network from port 12 to port 16
R16_12 nt_p_12 nt_c_16 337.83161479823934
X1507 nt_p_12 nt_c_16 rl_admittance res=158.59336007919467 ind=1.3684637459348558e-05
X1508 nt_n_12 nt_c_16 rl_admittance res=113.94021614950532 ind=4.355324314311421e-05
X1509 nt_n_12 nt_c_16 rl_admittance res=1540.374077463362 ind=0.0012931056943796797
X1510 nt_p_12 nt_c_16 rl_admittance res=343.1773783586659 ind=0.011664746367693282
X1511 nt_p_12 nt_c_16 rl_admittance res=54.55343221848019 ind=0.211789794889202
X1512 nt_n_12 nt_c_16 rl_admittance res=47.428371290047835 ind=0.015797489126330232
* Transfer network from port 13 to port 16
R16_13 nt_p_13 nt_c_16 535.212776405815
X1513 nt_n_13 nt_c_16 rl_admittance res=249.33372498677087 ind=2.1514404078008373e-05
X1514 nt_n_13 nt_c_16 rl_admittance res=1970.3276077262517 ind=0.0007531507335240787
X1515 nt_p_13 nt_c_16 rl_admittance res=359.65985362156135 ind=0.00030192549430829084
X1516 nt_n_13 nt_c_16 rl_admittance res=1086.5360368449963 ind=0.036931826187882745
X1517 nt_p_13 nt_c_16 rl_admittance res=90.05566603968427 ind=0.3496181681616395
X1518 nt_n_13 nt_c_16 rl_admittance res=96.95197713181597 ind=0.032292861063046116
* Transfer network from port 14 to port 16
R16_14 nt_p_14 nt_c_16 250.09738284267223
X1519 nt_n_14 nt_c_16 rl_admittance res=53.972810066263136 ind=4.657183239262131e-06
X1520 nt_p_14 nt_c_16 rl_admittance res=108.69283311928531 ind=4.1547449607666236e-05
X1521 nt_p_14 nt_c_16 rl_admittance res=189.27715745827706 ind=0.00015889346211820998
X1522 nt_p_14 nt_c_16 rl_admittance res=644.9958391341908 ind=0.02192368537722948
X1523 nt_p_14 nt_c_16 rl_admittance res=26.84927347053441 ind=0.10423546035518338
X1524 nt_n_14 nt_c_16 rl_admittance res=25.806762081902054 ind=0.00859574200601287
* Transfer network from port 15 to port 16
R16_15 nt_n_15 nt_c_16 4009.6200760746265
X1525 nt_n_15 nt_c_16 rl_admittance res=3634.324062238804 ind=0.0003135970331714376
X1526 nt_p_15 nt_c_16 rl_admittance res=1436.987556741172 ind=0.0005492833923560151
X1527 nt_n_15 nt_c_16 rl_admittance res=3462.986099437299 ind=0.0029070906283454752
X1528 nt_p_15 nt_c_16 rl_admittance res=569.7970888164072 ind=0.01936764758179042
X1529 nt_p_15 nt_c_16 rl_admittance res=76.69722862878723 ind=0.29775743998667176
X1530 nt_n_15 nt_c_16 rl_admittance res=68.13905848383385 ind=0.02269582543524149
* Transfer network from port 16 to port 16
R16_16 nt_p_16 nt_c_16 47.433503403105014
X1531 nt_n_16 nt_c_16 rl_admittance res=0.9242573367703678 ind=7.975193013458812e-08
X1532 nt_p_16 nt_c_16 rl_admittance res=13.692017351695982 ind=5.23372502695347e-06
X1533 nt_n_16 nt_c_16 rl_admittance res=91.08066509944268 ind=7.645995113208417e-05
X1534 nt_n_16 nt_c_16 rl_admittance res=600.1058762220235 ind=0.020397856272962808
X1535 nt_p_16 nt_c_16 rl_admittance res=523.0185859371131 ind=2.030486342183579
X1536 nt_n_16 nt_c_16 rl_admittance res=2304.2976792479694 ind=0.767517765034159
.ENDS s_equivalent

.SUBCKT rcl_vccs_admittance n_pos n_neg res=1e3 cap=1e-9 ind=100e-12 gm=1e-3
L1 n_pos 1 {ind}
C1 1 2 {cap}
R1 2 n_neg {res}
G1 n_pos n_neg 1 2 {gm}
.ENDS rcl_vccs_admittance

.SUBCKT rl_admittance n_pos n_neg res=1e3 ind=100e-12
L1 n_pos 1 {ind}
R1 1 n_neg {res}
.ENDS rl_admittance

